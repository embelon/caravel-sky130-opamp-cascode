magic
tech sky130A
magscale 1 2
timestamp 1698658818
<< nwell >>
rect 1066 114501 114670 115067
rect 1066 113413 114670 113979
rect 1066 112325 114670 112891
rect 1066 111237 114670 111803
rect 1066 110149 114670 110715
rect 1066 109061 114670 109627
rect 1066 107973 114670 108539
rect 1066 106885 114670 107451
rect 1066 105797 114670 106363
rect 1066 104709 114670 105275
rect 1066 103621 114670 104187
rect 1066 102533 114670 103099
rect 1066 101445 114670 102011
rect 1066 100357 114670 100923
rect 1066 99269 114670 99835
rect 1066 98181 114670 98747
rect 1066 97093 114670 97659
rect 1066 96005 114670 96571
rect 1066 94917 114670 95483
rect 1066 93829 114670 94395
rect 1066 92741 114670 93307
rect 1066 91653 114670 92219
rect 1066 90565 114670 91131
rect 1066 89477 114670 90043
rect 1066 88389 114670 88955
rect 1066 87301 114670 87867
rect 1066 86213 114670 86779
rect 1066 85125 114670 85691
rect 1066 84037 114670 84603
rect 1066 82949 114670 83515
rect 1066 81861 114670 82427
rect 1066 80773 114670 81339
rect 1066 79685 114670 80251
rect 1066 78597 114670 79163
rect 1066 77509 114670 78075
rect 1066 76421 114670 76987
rect 1066 75333 114670 75899
rect 1066 74245 114670 74811
rect 1066 73157 114670 73723
rect 1066 72069 114670 72635
rect 1066 70981 114670 71547
rect 1066 69893 114670 70459
rect 1066 68805 114670 69371
rect 1066 67717 114670 68283
rect 1066 66629 114670 67195
rect 1066 65541 114670 66107
rect 1066 64453 114670 65019
rect 1066 63365 114670 63931
rect 1066 62277 114670 62843
rect 1066 61189 114670 61755
rect 1066 60101 114670 60667
rect 1066 59013 114670 59579
rect 1066 57925 114670 58491
rect 1066 56837 114670 57403
rect 1066 55749 114670 56315
rect 1066 54661 114670 55227
rect 1066 53573 114670 54139
rect 1066 52485 114670 53051
rect 1066 51397 114670 51963
rect 1066 50309 114670 50875
rect 1066 49221 114670 49787
rect 1066 48133 114670 48699
rect 1066 47045 114670 47611
rect 1066 45957 114670 46523
rect 1066 44869 114670 45435
rect 1066 43781 114670 44347
rect 1066 42693 114670 43259
rect 1066 41605 114670 42171
rect 1066 40517 114670 41083
rect 1066 39429 114670 39995
rect 1066 38341 114670 38907
rect 1066 37253 114670 37819
rect 1066 36165 114670 36731
rect 1066 35077 114670 35643
rect 1066 33989 114670 34555
rect 1066 32901 114670 33467
rect 1066 31813 114670 32379
rect 1066 30725 114670 31291
rect 1066 29637 114670 30203
rect 1066 28549 114670 29115
rect 1066 27461 114670 28027
rect 1066 26373 114670 26939
rect 1066 25285 114670 25851
rect 1066 24197 114670 24763
rect 1066 23109 114670 23675
rect 1066 22021 114670 22587
rect 1066 20933 114670 21499
rect 1066 19845 114670 20411
rect 1066 18757 114670 19323
rect 1066 17669 114670 18235
rect 1066 16581 114670 17147
rect 1066 15493 114670 16059
rect 1066 14405 114670 14971
rect 1066 13317 114670 13883
rect 1066 12229 114670 12795
rect 1066 11141 114670 11707
rect 1066 10053 114670 10619
rect 1066 8965 114670 9531
rect 1066 7877 114670 8443
rect 1066 6789 114670 7355
rect 1066 5701 114670 6267
rect 1066 4613 114670 5179
rect 1066 3525 114670 4091
rect 1066 2437 114670 3003
<< obsli1 >>
rect 1104 2159 114632 115345
<< obsm1 >>
rect 1104 2128 114692 115456
<< metal2 >>
rect 1582 117118 1638 117918
rect 3974 117118 4030 117918
rect 6366 117118 6422 117918
rect 8758 117118 8814 117918
rect 11150 117118 11206 117918
rect 13542 117118 13598 117918
rect 15934 117118 15990 117918
rect 18326 117118 18382 117918
rect 20718 117118 20774 117918
rect 23110 117118 23166 117918
rect 25502 117118 25558 117918
rect 27894 117118 27950 117918
rect 30286 117118 30342 117918
rect 32678 117118 32734 117918
rect 35070 117118 35126 117918
rect 37462 117118 37518 117918
rect 39854 117118 39910 117918
rect 42246 117118 42302 117918
rect 44638 117118 44694 117918
rect 47030 117118 47086 117918
rect 49422 117118 49478 117918
rect 51814 117118 51870 117918
rect 54206 117118 54262 117918
rect 56598 117118 56654 117918
rect 58990 117118 59046 117918
rect 61382 117118 61438 117918
rect 63774 117118 63830 117918
rect 66166 117118 66222 117918
rect 68558 117118 68614 117918
rect 70950 117118 71006 117918
rect 73342 117118 73398 117918
rect 75734 117118 75790 117918
rect 78126 117118 78182 117918
rect 80518 117118 80574 117918
rect 82910 117118 82966 117918
rect 85302 117118 85358 117918
rect 87694 117118 87750 117918
rect 90086 117118 90142 117918
rect 92478 117118 92534 117918
rect 94870 117118 94926 117918
rect 97262 117118 97318 117918
rect 99654 117118 99710 117918
rect 102046 117118 102102 117918
rect 104438 117118 104494 117918
rect 106830 117118 106886 117918
rect 109222 117118 109278 117918
rect 111614 117118 111670 117918
rect 114006 117118 114062 117918
rect 1674 0 1730 800
rect 4710 0 4766 800
rect 7746 0 7802 800
rect 10782 0 10838 800
rect 13818 0 13874 800
rect 16854 0 16910 800
rect 19890 0 19946 800
rect 22926 0 22982 800
rect 25962 0 26018 800
rect 28998 0 29054 800
rect 32034 0 32090 800
rect 35070 0 35126 800
rect 38106 0 38162 800
rect 41142 0 41198 800
rect 44178 0 44234 800
rect 47214 0 47270 800
rect 50250 0 50306 800
rect 53286 0 53342 800
rect 56322 0 56378 800
rect 59358 0 59414 800
rect 62394 0 62450 800
rect 65430 0 65486 800
rect 68466 0 68522 800
rect 71502 0 71558 800
rect 74538 0 74594 800
rect 77574 0 77630 800
rect 80610 0 80666 800
rect 83646 0 83702 800
rect 86682 0 86738 800
rect 89718 0 89774 800
rect 92754 0 92810 800
rect 95790 0 95846 800
rect 98826 0 98882 800
rect 101862 0 101918 800
rect 104898 0 104954 800
rect 107934 0 107990 800
rect 110970 0 111026 800
rect 114006 0 114062 800
<< obsm2 >>
rect 1694 117062 3918 117118
rect 4086 117062 6310 117118
rect 6478 117062 8702 117118
rect 8870 117062 11094 117118
rect 11262 117062 13486 117118
rect 13654 117062 15878 117118
rect 16046 117062 18270 117118
rect 18438 117062 20662 117118
rect 20830 117062 23054 117118
rect 23222 117062 25446 117118
rect 25614 117062 27838 117118
rect 28006 117062 30230 117118
rect 30398 117062 32622 117118
rect 32790 117062 35014 117118
rect 35182 117062 37406 117118
rect 37574 117062 39798 117118
rect 39966 117062 42190 117118
rect 42358 117062 44582 117118
rect 44750 117062 46974 117118
rect 47142 117062 49366 117118
rect 49534 117062 51758 117118
rect 51926 117062 54150 117118
rect 54318 117062 56542 117118
rect 56710 117062 58934 117118
rect 59102 117062 61326 117118
rect 61494 117062 63718 117118
rect 63886 117062 66110 117118
rect 66278 117062 68502 117118
rect 68670 117062 70894 117118
rect 71062 117062 73286 117118
rect 73454 117062 75678 117118
rect 75846 117062 78070 117118
rect 78238 117062 80462 117118
rect 80630 117062 82854 117118
rect 83022 117062 85246 117118
rect 85414 117062 87638 117118
rect 87806 117062 90030 117118
rect 90198 117062 92422 117118
rect 92590 117062 94814 117118
rect 94982 117062 97206 117118
rect 97374 117062 99598 117118
rect 99766 117062 101990 117118
rect 102158 117062 104382 117118
rect 104550 117062 106774 117118
rect 106942 117062 109166 117118
rect 109334 117062 111558 117118
rect 111726 117062 113950 117118
rect 114118 117062 114336 117118
rect 1584 856 114336 117062
rect 1584 800 1618 856
rect 1786 800 4654 856
rect 4822 800 7690 856
rect 7858 800 10726 856
rect 10894 800 13762 856
rect 13930 800 16798 856
rect 16966 800 19834 856
rect 20002 800 22870 856
rect 23038 800 25906 856
rect 26074 800 28942 856
rect 29110 800 31978 856
rect 32146 800 35014 856
rect 35182 800 38050 856
rect 38218 800 41086 856
rect 41254 800 44122 856
rect 44290 800 47158 856
rect 47326 800 50194 856
rect 50362 800 53230 856
rect 53398 800 56266 856
rect 56434 800 59302 856
rect 59470 800 62338 856
rect 62506 800 65374 856
rect 65542 800 68410 856
rect 68578 800 71446 856
rect 71614 800 74482 856
rect 74650 800 77518 856
rect 77686 800 80554 856
rect 80722 800 83590 856
rect 83758 800 86626 856
rect 86794 800 89662 856
rect 89830 800 92698 856
rect 92866 800 95734 856
rect 95902 800 98770 856
rect 98938 800 101806 856
rect 101974 800 104842 856
rect 105010 800 107878 856
rect 108046 800 110914 856
rect 111082 800 113950 856
rect 114118 800 114336 856
<< metal3 >>
rect 114974 115744 115774 115864
rect 114974 112752 115774 112872
rect 114974 109760 115774 109880
rect 114974 106768 115774 106888
rect 114974 103776 115774 103896
rect 114974 100784 115774 100904
rect 114974 97792 115774 97912
rect 114974 94800 115774 94920
rect 114974 91808 115774 91928
rect 114974 88816 115774 88936
rect 114974 85824 115774 85944
rect 114974 82832 115774 82952
rect 114974 79840 115774 79960
rect 114974 76848 115774 76968
rect 114974 73856 115774 73976
rect 114974 70864 115774 70984
rect 114974 67872 115774 67992
rect 114974 64880 115774 65000
rect 114974 61888 115774 62008
rect 114974 58896 115774 59016
rect 114974 55904 115774 56024
rect 114974 52912 115774 53032
rect 114974 49920 115774 50040
rect 114974 46928 115774 47048
rect 114974 43936 115774 44056
rect 114974 40944 115774 41064
rect 114974 37952 115774 38072
rect 114974 34960 115774 35080
rect 114974 31968 115774 32088
rect 114974 28976 115774 29096
rect 114974 25984 115774 26104
rect 114974 22992 115774 23112
rect 114974 20000 115774 20120
rect 114974 17008 115774 17128
rect 114974 14016 115774 14136
rect 114974 11024 115774 11144
rect 114974 8032 115774 8152
rect 114974 5040 115774 5160
rect 114974 2048 115774 2168
<< obsm3 >>
rect 4210 115664 114894 115837
rect 4210 112952 114974 115664
rect 4210 112672 114894 112952
rect 4210 109960 114974 112672
rect 4210 109680 114894 109960
rect 4210 106968 114974 109680
rect 4210 106688 114894 106968
rect 4210 103976 114974 106688
rect 4210 103696 114894 103976
rect 4210 100984 114974 103696
rect 4210 100704 114894 100984
rect 4210 97992 114974 100704
rect 4210 97712 114894 97992
rect 4210 95000 114974 97712
rect 4210 94720 114894 95000
rect 4210 92008 114974 94720
rect 4210 91728 114894 92008
rect 4210 89016 114974 91728
rect 4210 88736 114894 89016
rect 4210 86024 114974 88736
rect 4210 85744 114894 86024
rect 4210 83032 114974 85744
rect 4210 82752 114894 83032
rect 4210 80040 114974 82752
rect 4210 79760 114894 80040
rect 4210 77048 114974 79760
rect 4210 76768 114894 77048
rect 4210 74056 114974 76768
rect 4210 73776 114894 74056
rect 4210 71064 114974 73776
rect 4210 70784 114894 71064
rect 4210 68072 114974 70784
rect 4210 67792 114894 68072
rect 4210 65080 114974 67792
rect 4210 64800 114894 65080
rect 4210 62088 114974 64800
rect 4210 61808 114894 62088
rect 4210 59096 114974 61808
rect 4210 58816 114894 59096
rect 4210 56104 114974 58816
rect 4210 55824 114894 56104
rect 4210 53112 114974 55824
rect 4210 52832 114894 53112
rect 4210 50120 114974 52832
rect 4210 49840 114894 50120
rect 4210 47128 114974 49840
rect 4210 46848 114894 47128
rect 4210 44136 114974 46848
rect 4210 43856 114894 44136
rect 4210 41144 114974 43856
rect 4210 40864 114894 41144
rect 4210 38152 114974 40864
rect 4210 37872 114894 38152
rect 4210 35160 114974 37872
rect 4210 34880 114894 35160
rect 4210 32168 114974 34880
rect 4210 31888 114894 32168
rect 4210 29176 114974 31888
rect 4210 28896 114894 29176
rect 4210 26184 114974 28896
rect 4210 25904 114894 26184
rect 4210 23192 114974 25904
rect 4210 22912 114894 23192
rect 4210 20200 114974 22912
rect 4210 19920 114894 20200
rect 4210 17208 114974 19920
rect 4210 16928 114894 17208
rect 4210 14216 114974 16928
rect 4210 13936 114894 14216
rect 4210 11224 114974 13936
rect 4210 10944 114894 11224
rect 4210 8232 114974 10944
rect 4210 7952 114894 8232
rect 4210 5240 114974 7952
rect 4210 4960 114894 5240
rect 4210 2248 114974 4960
rect 4210 1968 114894 2248
rect 4210 1939 114974 1968
<< metal4 >>
rect 4208 2128 4528 115376
rect 19568 2128 19888 115376
rect 34928 2128 35248 115376
rect 50288 2128 50608 115376
rect 65648 2128 65968 115376
rect 81008 2128 81328 115376
rect 96368 2128 96688 115376
rect 111728 2128 112048 115376
<< obsm4 >>
rect 15699 2048 19488 113389
rect 19968 2048 34848 113389
rect 35328 2048 50208 113389
rect 50688 2048 65568 113389
rect 66048 2048 80928 113389
rect 81408 2048 96288 113389
rect 96768 2048 98565 113389
rect 15699 1939 98565 2048
<< labels >>
rlabel metal3 s 114974 2048 115774 2168 6 i_clk
port 1 nsew signal input
rlabel metal3 s 114974 70864 115774 70984 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 114974 49920 115774 50040 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 114974 14016 115774 14136 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 114974 17008 115774 17128 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 114974 20000 115774 20120 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 114974 22992 115774 23112 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 114974 25984 115774 26104 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 114974 28976 115774 29096 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 114974 31968 115774 32088 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 114974 34960 115774 35080 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 114974 37952 115774 38072 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 114974 40944 115774 41064 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 114974 43936 115774 44056 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 114974 46928 115774 47048 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 114974 52912 115774 53032 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 114974 55904 115774 56024 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 114974 58896 115774 59016 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 114974 61888 115774 62008 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 114974 64880 115774 65000 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 114974 67872 115774 67992 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 114974 73856 115774 73976 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 114974 76848 115774 76968 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 114974 79840 115774 79960 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 114974 82832 115774 82952 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 114974 85824 115774 85944 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 114974 88816 115774 88936 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 114974 91808 115774 91928 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 114974 94800 115774 94920 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 114974 97792 115774 97912 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 114974 100784 115774 100904 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 114974 103776 115774 103896 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 114974 106768 115774 106888 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 114974 109760 115774 109880 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 114974 112752 115774 112872 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 114974 115744 115774 115864 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 114974 5040 115774 5160 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 114974 8032 115774 8152 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 114974 11024 115774 11144 6 i_reg_sclk
port 47 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 i_reset_lock_a
port 48 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 i_reset_lock_b
port 49 nsew signal input
rlabel metal2 s 8758 117118 8814 117918 6 i_tex_in[0]
port 50 nsew signal input
rlabel metal2 s 6366 117118 6422 117918 6 i_tex_in[1]
port 51 nsew signal input
rlabel metal2 s 3974 117118 4030 117918 6 i_tex_in[2]
port 52 nsew signal input
rlabel metal2 s 1582 117118 1638 117918 6 i_tex_in[3]
port 53 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 i_vec_csb
port 54 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 i_vec_mosi
port 55 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 i_vec_sclk
port 56 nsew signal input
rlabel metal2 s 23110 117118 23166 117918 6 o_gpout[0]
port 57 nsew signal output
rlabel metal2 s 20718 117118 20774 117918 6 o_gpout[1]
port 58 nsew signal output
rlabel metal2 s 18326 117118 18382 117918 6 o_gpout[2]
port 59 nsew signal output
rlabel metal2 s 15934 117118 15990 117918 6 o_gpout[3]
port 60 nsew signal output
rlabel metal2 s 13542 117118 13598 117918 6 o_gpout[4]
port 61 nsew signal output
rlabel metal2 s 11150 117118 11206 117918 6 o_gpout[5]
port 62 nsew signal output
rlabel metal2 s 37462 117118 37518 117918 6 o_hsync
port 63 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 o_reset
port 64 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 o_rgb[0]
port 65 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 o_rgb[10]
port 66 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 o_rgb[11]
port 67 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 o_rgb[12]
port 68 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 o_rgb[13]
port 69 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 o_rgb[14]
port 70 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 o_rgb[15]
port 71 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 o_rgb[16]
port 72 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 o_rgb[17]
port 73 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 o_rgb[18]
port 74 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 o_rgb[19]
port 75 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 o_rgb[1]
port 76 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 o_rgb[20]
port 77 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 o_rgb[21]
port 78 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 o_rgb[22]
port 79 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 o_rgb[23]
port 80 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 o_rgb[2]
port 81 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 o_rgb[3]
port 82 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 o_rgb[4]
port 83 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 o_rgb[5]
port 84 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 o_rgb[6]
port 85 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 o_rgb[7]
port 86 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 o_rgb[8]
port 87 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 o_rgb[9]
port 88 nsew signal output
rlabel metal2 s 32678 117118 32734 117918 6 o_tex_csb
port 89 nsew signal output
rlabel metal2 s 30286 117118 30342 117918 6 o_tex_oeb0
port 90 nsew signal output
rlabel metal2 s 27894 117118 27950 117918 6 o_tex_out0
port 91 nsew signal output
rlabel metal2 s 25502 117118 25558 117918 6 o_tex_sclk
port 92 nsew signal output
rlabel metal2 s 35070 117118 35126 117918 6 o_vsync
port 93 nsew signal output
rlabel metal2 s 114006 117118 114062 117918 6 ones[0]
port 94 nsew signal output
rlabel metal2 s 90086 117118 90142 117918 6 ones[10]
port 95 nsew signal output
rlabel metal2 s 87694 117118 87750 117918 6 ones[11]
port 96 nsew signal output
rlabel metal2 s 85302 117118 85358 117918 6 ones[12]
port 97 nsew signal output
rlabel metal2 s 82910 117118 82966 117918 6 ones[13]
port 98 nsew signal output
rlabel metal2 s 80518 117118 80574 117918 6 ones[14]
port 99 nsew signal output
rlabel metal2 s 78126 117118 78182 117918 6 ones[15]
port 100 nsew signal output
rlabel metal2 s 111614 117118 111670 117918 6 ones[1]
port 101 nsew signal output
rlabel metal2 s 109222 117118 109278 117918 6 ones[2]
port 102 nsew signal output
rlabel metal2 s 106830 117118 106886 117918 6 ones[3]
port 103 nsew signal output
rlabel metal2 s 104438 117118 104494 117918 6 ones[4]
port 104 nsew signal output
rlabel metal2 s 102046 117118 102102 117918 6 ones[5]
port 105 nsew signal output
rlabel metal2 s 99654 117118 99710 117918 6 ones[6]
port 106 nsew signal output
rlabel metal2 s 97262 117118 97318 117918 6 ones[7]
port 107 nsew signal output
rlabel metal2 s 94870 117118 94926 117918 6 ones[8]
port 108 nsew signal output
rlabel metal2 s 92478 117118 92534 117918 6 ones[9]
port 109 nsew signal output
rlabel metal4 s 4208 2128 4528 115376 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 115376 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 115376 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 115376 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 115376 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 115376 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 115376 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 115376 6 vssd1
port 111 nsew ground bidirectional
rlabel metal2 s 75734 117118 75790 117918 6 zeros[0]
port 112 nsew signal output
rlabel metal2 s 51814 117118 51870 117918 6 zeros[10]
port 113 nsew signal output
rlabel metal2 s 49422 117118 49478 117918 6 zeros[11]
port 114 nsew signal output
rlabel metal2 s 47030 117118 47086 117918 6 zeros[12]
port 115 nsew signal output
rlabel metal2 s 44638 117118 44694 117918 6 zeros[13]
port 116 nsew signal output
rlabel metal2 s 42246 117118 42302 117918 6 zeros[14]
port 117 nsew signal output
rlabel metal2 s 39854 117118 39910 117918 6 zeros[15]
port 118 nsew signal output
rlabel metal2 s 73342 117118 73398 117918 6 zeros[1]
port 119 nsew signal output
rlabel metal2 s 70950 117118 71006 117918 6 zeros[2]
port 120 nsew signal output
rlabel metal2 s 68558 117118 68614 117918 6 zeros[3]
port 121 nsew signal output
rlabel metal2 s 66166 117118 66222 117918 6 zeros[4]
port 122 nsew signal output
rlabel metal2 s 63774 117118 63830 117918 6 zeros[5]
port 123 nsew signal output
rlabel metal2 s 61382 117118 61438 117918 6 zeros[6]
port 124 nsew signal output
rlabel metal2 s 58990 117118 59046 117918 6 zeros[7]
port 125 nsew signal output
rlabel metal2 s 56598 117118 56654 117918 6 zeros[8]
port 126 nsew signal output
rlabel metal2 s 54206 117118 54262 117918 6 zeros[9]
port 127 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 115774 117918
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32187136
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_10_30_20_05/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1535530
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 587.570 BY 598.290 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 12.960 587.570 13.560 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 355.680 587.570 356.280 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 255.720 587.570 256.320 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 84.360 587.570 84.960 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 98.640 587.570 99.240 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 112.920 587.570 113.520 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 127.200 587.570 127.800 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 141.480 587.570 142.080 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 155.760 587.570 156.360 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 170.040 587.570 170.640 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 184.320 587.570 184.920 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 198.600 587.570 199.200 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 212.880 587.570 213.480 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 227.160 587.570 227.760 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 241.440 587.570 242.040 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 270.000 587.570 270.600 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 284.280 587.570 284.880 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 298.560 587.570 299.160 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 312.840 587.570 313.440 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 327.120 587.570 327.720 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 341.400 587.570 342.000 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 369.960 587.570 370.560 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 384.240 587.570 384.840 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 398.520 587.570 399.120 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 412.800 587.570 413.400 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 427.080 587.570 427.680 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 441.360 587.570 441.960 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 455.640 587.570 456.240 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 469.920 587.570 470.520 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 484.200 587.570 484.800 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 498.480 587.570 499.080 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 512.760 587.570 513.360 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 527.040 587.570 527.640 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 541.320 587.570 541.920 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 555.600 587.570 556.200 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 569.880 587.570 570.480 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 27.240 587.570 27.840 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 41.520 587.570 42.120 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 55.800 587.570 56.400 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 70.080 587.570 70.680 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.570 584.160 587.570 584.760 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 594.290 6.810 598.290 ;
    END
  END i_spare_1
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 594.290 54.650 598.290 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 594.290 42.690 598.290 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 594.290 30.730 598.290 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 594.290 18.770 598.290 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 594.290 126.410 598.290 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 594.290 114.450 598.290 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 594.290 102.490 598.290 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 594.290 90.530 598.290 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 594.290 78.570 598.290 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 594.290 66.610 598.290 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 594.290 198.170 598.290 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 594.290 174.250 598.290 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 594.290 162.290 598.290 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 594.290 150.330 598.290 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 594.290 138.370 598.290 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 594.290 186.210 598.290 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 594.290 580.890 598.290 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 594.290 461.290 598.290 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 594.290 449.330 598.290 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 594.290 437.370 598.290 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 594.290 425.410 598.290 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 594.290 413.450 598.290 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 594.290 401.490 598.290 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 594.290 568.930 598.290 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 594.290 556.970 598.290 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 594.290 545.010 598.290 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 594.290 533.050 598.290 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 594.290 521.090 598.290 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 594.290 509.130 598.290 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 594.290 497.170 598.290 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 594.290 485.210 598.290 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 594.290 473.250 598.290 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 585.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 585.040 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 594.290 389.530 598.290 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 594.290 269.930 598.290 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 594.290 257.970 598.290 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 594.290 246.010 598.290 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 594.290 234.050 598.290 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 594.290 222.090 598.290 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 594.290 210.130 598.290 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 594.290 377.570 598.290 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 594.290 365.610 598.290 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 594.290 353.650 598.290 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 594.290 341.690 598.290 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 594.290 329.730 598.290 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 594.290 317.770 598.290 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 594.290 305.810 598.290 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 594.290 293.850 598.290 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 594.290 281.890 598.290 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 582.090 584.990 ;
        RECT 5.330 577.945 582.090 580.775 ;
        RECT 5.330 572.505 582.090 575.335 ;
        RECT 5.330 567.065 582.090 569.895 ;
        RECT 5.330 561.625 582.090 564.455 ;
        RECT 5.330 556.185 582.090 559.015 ;
        RECT 5.330 550.745 582.090 553.575 ;
        RECT 5.330 545.305 582.090 548.135 ;
        RECT 5.330 539.865 582.090 542.695 ;
        RECT 5.330 534.425 582.090 537.255 ;
        RECT 5.330 528.985 582.090 531.815 ;
        RECT 5.330 523.545 582.090 526.375 ;
        RECT 5.330 518.105 582.090 520.935 ;
        RECT 5.330 512.665 582.090 515.495 ;
        RECT 5.330 507.225 582.090 510.055 ;
        RECT 5.330 501.785 582.090 504.615 ;
        RECT 5.330 496.345 582.090 499.175 ;
        RECT 5.330 490.905 582.090 493.735 ;
        RECT 5.330 485.465 582.090 488.295 ;
        RECT 5.330 480.025 582.090 482.855 ;
        RECT 5.330 474.585 582.090 477.415 ;
        RECT 5.330 469.145 582.090 471.975 ;
        RECT 5.330 463.705 582.090 466.535 ;
        RECT 5.330 458.265 582.090 461.095 ;
        RECT 5.330 452.825 582.090 455.655 ;
        RECT 5.330 447.385 582.090 450.215 ;
        RECT 5.330 441.945 582.090 444.775 ;
        RECT 5.330 436.505 582.090 439.335 ;
        RECT 5.330 431.065 582.090 433.895 ;
        RECT 5.330 425.625 582.090 428.455 ;
        RECT 5.330 420.185 582.090 423.015 ;
        RECT 5.330 414.745 582.090 417.575 ;
        RECT 5.330 409.305 582.090 412.135 ;
        RECT 5.330 403.865 582.090 406.695 ;
        RECT 5.330 398.425 582.090 401.255 ;
        RECT 5.330 392.985 582.090 395.815 ;
        RECT 5.330 387.545 582.090 390.375 ;
        RECT 5.330 382.105 582.090 384.935 ;
        RECT 5.330 376.665 582.090 379.495 ;
        RECT 5.330 371.225 582.090 374.055 ;
        RECT 5.330 365.785 582.090 368.615 ;
        RECT 5.330 360.345 582.090 363.175 ;
        RECT 5.330 354.905 582.090 357.735 ;
        RECT 5.330 349.465 582.090 352.295 ;
        RECT 5.330 344.025 582.090 346.855 ;
        RECT 5.330 338.585 582.090 341.415 ;
        RECT 5.330 333.145 582.090 335.975 ;
        RECT 5.330 327.705 582.090 330.535 ;
        RECT 5.330 322.265 582.090 325.095 ;
        RECT 5.330 316.825 582.090 319.655 ;
        RECT 5.330 311.385 582.090 314.215 ;
        RECT 5.330 305.945 582.090 308.775 ;
        RECT 5.330 300.505 582.090 303.335 ;
        RECT 5.330 295.065 582.090 297.895 ;
        RECT 5.330 289.625 582.090 292.455 ;
        RECT 5.330 284.185 582.090 287.015 ;
        RECT 5.330 278.745 582.090 281.575 ;
        RECT 5.330 273.305 582.090 276.135 ;
        RECT 5.330 267.865 582.090 270.695 ;
        RECT 5.330 262.425 582.090 265.255 ;
        RECT 5.330 256.985 582.090 259.815 ;
        RECT 5.330 251.545 582.090 254.375 ;
        RECT 5.330 246.105 582.090 248.935 ;
        RECT 5.330 240.665 582.090 243.495 ;
        RECT 5.330 235.225 582.090 238.055 ;
        RECT 5.330 229.785 582.090 232.615 ;
        RECT 5.330 224.345 582.090 227.175 ;
        RECT 5.330 218.905 582.090 221.735 ;
        RECT 5.330 213.465 582.090 216.295 ;
        RECT 5.330 208.025 582.090 210.855 ;
        RECT 5.330 202.585 582.090 205.415 ;
        RECT 5.330 197.145 582.090 199.975 ;
        RECT 5.330 191.705 582.090 194.535 ;
        RECT 5.330 186.265 582.090 189.095 ;
        RECT 5.330 180.825 582.090 183.655 ;
        RECT 5.330 175.385 582.090 178.215 ;
        RECT 5.330 169.945 582.090 172.775 ;
        RECT 5.330 164.505 582.090 167.335 ;
        RECT 5.330 159.065 582.090 161.895 ;
        RECT 5.330 153.625 582.090 156.455 ;
        RECT 5.330 148.185 582.090 151.015 ;
        RECT 5.330 142.745 582.090 145.575 ;
        RECT 5.330 137.305 582.090 140.135 ;
        RECT 5.330 131.865 582.090 134.695 ;
        RECT 5.330 126.425 582.090 129.255 ;
        RECT 5.330 120.985 582.090 123.815 ;
        RECT 5.330 115.545 582.090 118.375 ;
        RECT 5.330 110.105 582.090 112.935 ;
        RECT 5.330 104.665 582.090 107.495 ;
        RECT 5.330 99.225 582.090 102.055 ;
        RECT 5.330 93.785 582.090 96.615 ;
        RECT 5.330 88.345 582.090 91.175 ;
        RECT 5.330 82.905 582.090 85.735 ;
        RECT 5.330 77.465 582.090 80.295 ;
        RECT 5.330 72.025 582.090 74.855 ;
        RECT 5.330 66.585 582.090 69.415 ;
        RECT 5.330 61.145 582.090 63.975 ;
        RECT 5.330 55.705 582.090 58.535 ;
        RECT 5.330 50.265 582.090 53.095 ;
        RECT 5.330 44.825 582.090 47.655 ;
        RECT 5.330 39.385 582.090 42.215 ;
        RECT 5.330 33.945 582.090 36.775 ;
        RECT 5.330 28.505 582.090 31.335 ;
        RECT 5.330 23.065 582.090 25.895 ;
        RECT 5.330 17.625 582.090 20.455 ;
        RECT 5.330 12.185 582.090 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 581.900 584.885 ;
      LAYER met1 ;
        RECT 5.520 9.220 581.900 585.040 ;
      LAYER met2 ;
        RECT 7.920 594.010 18.210 594.290 ;
        RECT 19.050 594.010 30.170 594.290 ;
        RECT 31.010 594.010 42.130 594.290 ;
        RECT 42.970 594.010 54.090 594.290 ;
        RECT 54.930 594.010 66.050 594.290 ;
        RECT 66.890 594.010 78.010 594.290 ;
        RECT 78.850 594.010 89.970 594.290 ;
        RECT 90.810 594.010 101.930 594.290 ;
        RECT 102.770 594.010 113.890 594.290 ;
        RECT 114.730 594.010 125.850 594.290 ;
        RECT 126.690 594.010 137.810 594.290 ;
        RECT 138.650 594.010 149.770 594.290 ;
        RECT 150.610 594.010 161.730 594.290 ;
        RECT 162.570 594.010 173.690 594.290 ;
        RECT 174.530 594.010 185.650 594.290 ;
        RECT 186.490 594.010 197.610 594.290 ;
        RECT 198.450 594.010 209.570 594.290 ;
        RECT 210.410 594.010 221.530 594.290 ;
        RECT 222.370 594.010 233.490 594.290 ;
        RECT 234.330 594.010 245.450 594.290 ;
        RECT 246.290 594.010 257.410 594.290 ;
        RECT 258.250 594.010 269.370 594.290 ;
        RECT 270.210 594.010 281.330 594.290 ;
        RECT 282.170 594.010 293.290 594.290 ;
        RECT 294.130 594.010 305.250 594.290 ;
        RECT 306.090 594.010 317.210 594.290 ;
        RECT 318.050 594.010 329.170 594.290 ;
        RECT 330.010 594.010 341.130 594.290 ;
        RECT 341.970 594.010 353.090 594.290 ;
        RECT 353.930 594.010 365.050 594.290 ;
        RECT 365.890 594.010 377.010 594.290 ;
        RECT 377.850 594.010 388.970 594.290 ;
        RECT 389.810 594.010 400.930 594.290 ;
        RECT 401.770 594.010 412.890 594.290 ;
        RECT 413.730 594.010 424.850 594.290 ;
        RECT 425.690 594.010 436.810 594.290 ;
        RECT 437.650 594.010 448.770 594.290 ;
        RECT 449.610 594.010 460.730 594.290 ;
        RECT 461.570 594.010 472.690 594.290 ;
        RECT 473.530 594.010 484.650 594.290 ;
        RECT 485.490 594.010 496.610 594.290 ;
        RECT 497.450 594.010 508.570 594.290 ;
        RECT 509.410 594.010 520.530 594.290 ;
        RECT 521.370 594.010 532.490 594.290 ;
        RECT 533.330 594.010 544.450 594.290 ;
        RECT 545.290 594.010 556.410 594.290 ;
        RECT 557.250 594.010 568.370 594.290 ;
        RECT 569.210 594.010 580.330 594.290 ;
        RECT 7.920 4.280 580.880 594.010 ;
        RECT 7.920 3.670 12.230 4.280 ;
        RECT 13.070 3.670 27.410 4.280 ;
        RECT 28.250 3.670 42.590 4.280 ;
        RECT 43.430 3.670 57.770 4.280 ;
        RECT 58.610 3.670 72.950 4.280 ;
        RECT 73.790 3.670 88.130 4.280 ;
        RECT 88.970 3.670 103.310 4.280 ;
        RECT 104.150 3.670 118.490 4.280 ;
        RECT 119.330 3.670 133.670 4.280 ;
        RECT 134.510 3.670 148.850 4.280 ;
        RECT 149.690 3.670 164.030 4.280 ;
        RECT 164.870 3.670 179.210 4.280 ;
        RECT 180.050 3.670 194.390 4.280 ;
        RECT 195.230 3.670 209.570 4.280 ;
        RECT 210.410 3.670 224.750 4.280 ;
        RECT 225.590 3.670 239.930 4.280 ;
        RECT 240.770 3.670 255.110 4.280 ;
        RECT 255.950 3.670 270.290 4.280 ;
        RECT 271.130 3.670 285.470 4.280 ;
        RECT 286.310 3.670 300.650 4.280 ;
        RECT 301.490 3.670 315.830 4.280 ;
        RECT 316.670 3.670 331.010 4.280 ;
        RECT 331.850 3.670 346.190 4.280 ;
        RECT 347.030 3.670 361.370 4.280 ;
        RECT 362.210 3.670 376.550 4.280 ;
        RECT 377.390 3.670 391.730 4.280 ;
        RECT 392.570 3.670 406.910 4.280 ;
        RECT 407.750 3.670 422.090 4.280 ;
        RECT 422.930 3.670 437.270 4.280 ;
        RECT 438.110 3.670 452.450 4.280 ;
        RECT 453.290 3.670 467.630 4.280 ;
        RECT 468.470 3.670 482.810 4.280 ;
        RECT 483.650 3.670 497.990 4.280 ;
        RECT 498.830 3.670 513.170 4.280 ;
        RECT 514.010 3.670 528.350 4.280 ;
        RECT 529.190 3.670 543.530 4.280 ;
        RECT 544.370 3.670 558.710 4.280 ;
        RECT 559.550 3.670 573.890 4.280 ;
        RECT 574.730 3.670 580.880 4.280 ;
      LAYER met3 ;
        RECT 21.050 583.760 583.170 584.965 ;
        RECT 21.050 570.880 583.570 583.760 ;
        RECT 21.050 569.480 583.170 570.880 ;
        RECT 21.050 556.600 583.570 569.480 ;
        RECT 21.050 555.200 583.170 556.600 ;
        RECT 21.050 542.320 583.570 555.200 ;
        RECT 21.050 540.920 583.170 542.320 ;
        RECT 21.050 528.040 583.570 540.920 ;
        RECT 21.050 526.640 583.170 528.040 ;
        RECT 21.050 513.760 583.570 526.640 ;
        RECT 21.050 512.360 583.170 513.760 ;
        RECT 21.050 499.480 583.570 512.360 ;
        RECT 21.050 498.080 583.170 499.480 ;
        RECT 21.050 485.200 583.570 498.080 ;
        RECT 21.050 483.800 583.170 485.200 ;
        RECT 21.050 470.920 583.570 483.800 ;
        RECT 21.050 469.520 583.170 470.920 ;
        RECT 21.050 456.640 583.570 469.520 ;
        RECT 21.050 455.240 583.170 456.640 ;
        RECT 21.050 442.360 583.570 455.240 ;
        RECT 21.050 440.960 583.170 442.360 ;
        RECT 21.050 428.080 583.570 440.960 ;
        RECT 21.050 426.680 583.170 428.080 ;
        RECT 21.050 413.800 583.570 426.680 ;
        RECT 21.050 412.400 583.170 413.800 ;
        RECT 21.050 399.520 583.570 412.400 ;
        RECT 21.050 398.120 583.170 399.520 ;
        RECT 21.050 385.240 583.570 398.120 ;
        RECT 21.050 383.840 583.170 385.240 ;
        RECT 21.050 370.960 583.570 383.840 ;
        RECT 21.050 369.560 583.170 370.960 ;
        RECT 21.050 356.680 583.570 369.560 ;
        RECT 21.050 355.280 583.170 356.680 ;
        RECT 21.050 342.400 583.570 355.280 ;
        RECT 21.050 341.000 583.170 342.400 ;
        RECT 21.050 328.120 583.570 341.000 ;
        RECT 21.050 326.720 583.170 328.120 ;
        RECT 21.050 313.840 583.570 326.720 ;
        RECT 21.050 312.440 583.170 313.840 ;
        RECT 21.050 299.560 583.570 312.440 ;
        RECT 21.050 298.160 583.170 299.560 ;
        RECT 21.050 285.280 583.570 298.160 ;
        RECT 21.050 283.880 583.170 285.280 ;
        RECT 21.050 271.000 583.570 283.880 ;
        RECT 21.050 269.600 583.170 271.000 ;
        RECT 21.050 256.720 583.570 269.600 ;
        RECT 21.050 255.320 583.170 256.720 ;
        RECT 21.050 242.440 583.570 255.320 ;
        RECT 21.050 241.040 583.170 242.440 ;
        RECT 21.050 228.160 583.570 241.040 ;
        RECT 21.050 226.760 583.170 228.160 ;
        RECT 21.050 213.880 583.570 226.760 ;
        RECT 21.050 212.480 583.170 213.880 ;
        RECT 21.050 199.600 583.570 212.480 ;
        RECT 21.050 198.200 583.170 199.600 ;
        RECT 21.050 185.320 583.570 198.200 ;
        RECT 21.050 183.920 583.170 185.320 ;
        RECT 21.050 171.040 583.570 183.920 ;
        RECT 21.050 169.640 583.170 171.040 ;
        RECT 21.050 156.760 583.570 169.640 ;
        RECT 21.050 155.360 583.170 156.760 ;
        RECT 21.050 142.480 583.570 155.360 ;
        RECT 21.050 141.080 583.170 142.480 ;
        RECT 21.050 128.200 583.570 141.080 ;
        RECT 21.050 126.800 583.170 128.200 ;
        RECT 21.050 113.920 583.570 126.800 ;
        RECT 21.050 112.520 583.170 113.920 ;
        RECT 21.050 99.640 583.570 112.520 ;
        RECT 21.050 98.240 583.170 99.640 ;
        RECT 21.050 85.360 583.570 98.240 ;
        RECT 21.050 83.960 583.170 85.360 ;
        RECT 21.050 71.080 583.570 83.960 ;
        RECT 21.050 69.680 583.170 71.080 ;
        RECT 21.050 56.800 583.570 69.680 ;
        RECT 21.050 55.400 583.170 56.800 ;
        RECT 21.050 42.520 583.570 55.400 ;
        RECT 21.050 41.120 583.170 42.520 ;
        RECT 21.050 28.240 583.570 41.120 ;
        RECT 21.050 26.840 583.170 28.240 ;
        RECT 21.050 13.960 583.570 26.840 ;
        RECT 21.050 12.560 583.170 13.960 ;
        RECT 21.050 10.715 583.570 12.560 ;
      LAYER met4 ;
        RECT 131.855 12.415 174.240 583.265 ;
        RECT 176.640 12.415 251.040 583.265 ;
        RECT 253.440 12.415 327.840 583.265 ;
        RECT 330.240 12.415 404.640 583.265 ;
        RECT 407.040 12.415 481.440 583.265 ;
        RECT 483.840 12.415 558.240 583.265 ;
        RECT 560.640 12.415 576.545 583.265 ;
  END
END top_ew_algofoogle
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1698599793
<< nwell >>
rect 1066 44869 14850 45435
rect 1066 43781 14850 44347
rect 1066 42693 14850 43259
rect 1066 41605 14850 42171
rect 1066 40517 14850 41083
rect 1066 39429 14850 39995
rect 1066 38341 14850 38907
rect 1066 37253 14850 37819
rect 1066 36165 14850 36731
rect 1066 35077 14850 35643
rect 1066 33989 14850 34555
rect 1066 32901 14850 33467
rect 1066 31813 14850 32379
rect 1066 30725 14850 31291
rect 1066 29637 14850 30203
rect 1066 28549 14850 29115
rect 1066 27461 14850 28027
rect 1066 26373 14850 26939
rect 1066 25285 14850 25851
rect 1066 24197 14850 24763
rect 1066 23109 14850 23675
rect 1066 22021 14850 22587
rect 1066 20933 14850 21499
rect 1066 19845 14850 20411
rect 1066 18757 14850 19323
rect 1066 17669 14850 18235
rect 1066 16581 14850 17147
rect 1066 15493 14850 16059
rect 1066 14405 14850 14971
rect 1066 13317 14850 13883
rect 1066 12229 14850 12795
rect 1066 11141 14850 11707
rect 1066 10053 14850 10619
rect 1066 8965 14850 9531
rect 1066 7877 14850 8443
rect 1066 6789 14850 7355
rect 1066 5701 14850 6267
rect 1066 4613 14850 5179
rect 1066 3525 14850 4091
rect 1066 2437 14850 3003
<< obsli1 >>
rect 1104 2159 14812 45713
<< obsm1 >>
rect 1104 2128 14971 45744
<< obsm2 >>
rect 2663 2139 14965 45733
<< metal3 >>
rect 15200 44888 16000 45008
rect 15200 41080 16000 41200
rect 15200 37272 16000 37392
rect 15200 33464 16000 33584
rect 15200 29656 16000 29776
rect 15200 25848 16000 25968
rect 15200 22040 16000 22160
rect 15200 18232 16000 18352
rect 15200 14424 16000 14544
rect 15200 10616 16000 10736
rect 15200 6808 16000 6928
rect 15200 3000 16000 3120
<< obsm3 >>
rect 2659 45088 15200 45729
rect 2659 44808 15120 45088
rect 2659 41280 15200 44808
rect 2659 41000 15120 41280
rect 2659 37472 15200 41000
rect 2659 37192 15120 37472
rect 2659 33664 15200 37192
rect 2659 33384 15120 33664
rect 2659 29856 15200 33384
rect 2659 29576 15120 29856
rect 2659 26048 15200 29576
rect 2659 25768 15120 26048
rect 2659 22240 15200 25768
rect 2659 21960 15120 22240
rect 2659 18432 15200 21960
rect 2659 18152 15120 18432
rect 2659 14624 15200 18152
rect 2659 14344 15120 14624
rect 2659 10816 15200 14344
rect 2659 10536 15120 10816
rect 2659 7008 15200 10536
rect 2659 6728 15120 7008
rect 2659 3200 15200 6728
rect 2659 2920 15120 3200
rect 2659 2143 15200 2920
<< metal4 >>
rect 2657 2128 2977 45744
rect 4370 2128 4690 45744
rect 6084 2128 6404 45744
rect 7797 2128 8117 45744
rect 9511 2128 9831 45744
rect 11224 2128 11544 45744
rect 12938 2128 13258 45744
rect 14651 2128 14971 45744
<< labels >>
rlabel metal3 s 15200 6808 16000 6928 6 io_oeb[0]
port 1 nsew signal output
rlabel metal3 s 15200 14424 16000 14544 6 io_oeb[1]
port 2 nsew signal output
rlabel metal3 s 15200 22040 16000 22160 6 io_oeb[2]
port 3 nsew signal output
rlabel metal3 s 15200 29656 16000 29776 6 io_oeb[3]
port 4 nsew signal output
rlabel metal3 s 15200 37272 16000 37392 6 io_oeb[4]
port 5 nsew signal output
rlabel metal3 s 15200 44888 16000 45008 6 io_oeb[5]
port 6 nsew signal output
rlabel metal3 s 15200 3000 16000 3120 6 io_out[0]
port 7 nsew signal output
rlabel metal3 s 15200 10616 16000 10736 6 io_out[1]
port 8 nsew signal output
rlabel metal3 s 15200 18232 16000 18352 6 io_out[2]
port 9 nsew signal output
rlabel metal3 s 15200 25848 16000 25968 6 io_out[3]
port 10 nsew signal output
rlabel metal3 s 15200 33464 16000 33584 6 io_out[4]
port 11 nsew signal output
rlabel metal3 s 15200 41080 16000 41200 6 io_out[5]
port 12 nsew signal output
rlabel metal4 s 2657 2128 2977 45744 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 45744 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 45744 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 45744 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 45744 6 vssd1
port 14 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 45744 6 vssd1
port 14 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 45744 6 vssd1
port 14 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 45744 6 vssd1
port 14 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 48000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 487224
string GDS_FILE /home/zwierzak/projects/caravel_user_project/openlane/analog_io_control/runs/23_10_29_18_09/results/signoff/analog_io_control.magic.gds
string GDS_START 23768
<< end >>


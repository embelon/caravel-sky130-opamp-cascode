* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_la_invalid i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_outs_enb i_reg_sclk i_reset_lock_a i_reset_lock_b i_spare_0 i_spare_1 i_tex_in[0]
+ i_tex_in[1] i_tex_in[2] i_tex_in[3] i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1]
+ o_gpout[2] o_gpout[3] o_gpout[4] o_gpout[5] o_hsync o_reset o_rgb[0] o_rgb[10] o_rgb[11]
+ o_rgb[12] o_rgb[13] o_rgb[14] o_rgb[15] o_rgb[16] o_rgb[17] o_rgb[18] o_rgb[19]
+ o_rgb[1] o_rgb[20] o_rgb[21] o_rgb[22] o_rgb[23] o_rgb[2] o_rgb[3] o_rgb[4] o_rgb[5]
+ o_rgb[6] o_rgb[7] o_rgb[8] o_rgb[9] o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk o_vsync
+ ones[0] ones[10] ones[11] ones[12] ones[13] ones[14] ones[15] ones[1] ones[2] ones[3]
+ ones[4] ones[5] ones[6] ones[7] ones[8] ones[9] vccd1 vssd1 zeros[0] zeros[10] zeros[11]
+ zeros[12] zeros[13] zeros[14] zeros[15] zeros[1] zeros[2] zeros[3] zeros[4] zeros[5]
+ zeros[6] zeros[7] zeros[8] zeros[9]
XFILLER_67_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18869_ _03015_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20900_ clknet_leaf_53_i_clk _00489_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_21880_ net406 _01469_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
X_20831_ clknet_leaf_67_i_clk _00420_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_36_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20762_ rbzero.wall_tracer.rayAddendX\[-6\] _02606_ _02557_ _03948_ vssd1 vssd1 vccd1
+ vccd1 _01650_ sky130_fd_sc_hd__a22o_1
XFILLER_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20693_ _03903_ _03906_ _03904_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21314_ clknet_leaf_1_i_clk _00903_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21245_ clknet_leaf_26_i_clk _00834_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21176_ clknet_leaf_14_i_clk _00765_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20127_ rbzero.vga_sync.vsync _03718_ _03720_ _03703_ vssd1 vssd1 vccd1 vccd1 _01242_
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20058_ _03212_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__clkbuf_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _05088_ _05069_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__or2b_2
XFILLER_133_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12880_ _06008_ _06050_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__xor2_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ rbzero.row_render.texu\[3\] vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__inv_2
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _07719_ _07720_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__nand2_1
XFILLER_54_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _04918_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__clkbuf_8
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13501_ _06605_ _06659_ _06576_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__mux2_1
XFILLER_92_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10713_ _04147_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__clkbuf_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14481_ _07611_ _07609_ _07610_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__nand3_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ gpout0.hpos\[9\] _04863_ _04879_ _04881_ _04882_ vssd1 vssd1 vccd1 vccd1
+ _04883_ sky130_fd_sc_hd__o221a_1
X_16220_ _09307_ _09312_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__xor2_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13432_ _06571_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__clkbuf_4
X_10644_ rbzero.tex_r0\[14\] rbzero.tex_r0\[13\] _04110_ vssd1 vssd1 vccd1 vccd1 _04111_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16151_ _08616_ _09243_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__nor2_2
XFILLER_155_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10575_ _04074_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _06520_ _06532_ _06533_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a21bo_1
XFILLER_155_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ rbzero.side_hot _06358_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__nand2_1
X_12314_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _04907_ vssd1 vssd1 vccd1 vccd1 _05500_
+ sky130_fd_sc_hd__mux2_1
X_16082_ _08429_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__buf_2
XFILLER_170_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ _06408_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__xnor2_2
X_19910_ rbzero.debug_overlay.playerX\[-5\] _03569_ _03574_ _03302_ vssd1 vssd1 vccd1
+ vccd1 _01171_ sky130_fd_sc_hd__o211a_1
X_15033_ _08125_ _08129_ _08130_ _08085_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__o211a_1
X_12245_ rbzero.tex_g1\[58\] _04830_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__or2_1
XFILLER_107_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12176_ rbzero.tex_g0\[62\] _05002_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__and2_1
X_19841_ _03532_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11127_ _04364_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
X_16984_ _09717_ _10005_ vssd1 vssd1 vccd1 vccd1 _10006_ sky130_fd_sc_hd__xor2_4
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19772_ _03496_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15935_ _08368_ _08373_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__nor2_1
X_11058_ _04328_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
X_18723_ _02908_ _02911_ _02920_ _04434_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a211o_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20506__351 clknet_1_0__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__inv_2
XFILLER_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18654_ _02841_ _02854_ _02855_ _04433_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a31o_1
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _08296_ _08953_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__or2_1
XFILLER_149_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _01811_ _01812_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__nand2_1
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14817_ _07827_ _07858_ _07860_ _06580_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__a211o_1
X_18585_ rbzero.wall_tracer.rayAddendY\[-1\] _09744_ _02792_ _02534_ vssd1 vssd1 vccd1
+ vccd1 _02793_ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_120 vssd1 vssd1 vccd1 vccd1 ones[11] top_ew_algofoogle_120/LO sky130_fd_sc_hd__conb_1
X_15797_ _08888_ _08891_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__xnor2_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _01805_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__xnor2_1
X_14748_ _06665_ _07914_ _07915_ _06663_ _06602_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__o221a_1
XFILLER_205_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _09822_ _10379_ _10380_ _09812_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__o311a_1
X_14679_ _07837_ _07841_ _07848_ _07849_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__o31ai_4
XFILLER_33_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ _09507_ _09508_ vssd1 vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__nor2_1
X_19206_ rbzero.spi_registers.texadd2\[1\] _03208_ vssd1 vssd1 vccd1 vccd1 _03210_
+ sky130_fd_sc_hd__or2_1
X_17398_ _01689_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nand2_1
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19137_ rbzero.spi_registers.new_texadd\[0\]\[20\] _03140_ _03168_ _03169_ vssd1
+ vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__o211a_1
XFILLER_192_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16349_ _09305_ _09318_ _09440_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__a21o_1
XFILLER_146_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19068_ rbzero.spi_registers.new_mapd\[4\] _03120_ _03129_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00773_ sky130_fd_sc_hd__o211a_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20251__121 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__inv_2
XFILLER_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ _02304_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__nor2_1
XFILLER_156_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21030_ clknet_leaf_17_i_clk _00619_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21932_ net458 _01521_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21863_ net389 _01452_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20814_ clknet_leaf_62_i_clk _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_21794_ net320 _01383_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20745_ rbzero.traced_texVinit\[10\] _02606_ _02557_ _10258_ vssd1 vssd1 vccd1 vccd1
+ _01644_ sky130_fd_sc_hd__a22o_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20676_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__and2b_1
XFILLER_196_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12030_ rbzero.tex_r1\[28\] _05185_ _05195_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_
+ sky130_fd_sc_hd__a31o_1
XFILLER_151_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21228_ clknet_leaf_11_i_clk _00817_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21159_ clknet_leaf_12_i_clk _00748_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _07150_ _07151_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__nand2_1
XFILLER_59_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15720_ _08814_ _08696_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__or2_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12932_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__inv_2
XFILLER_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _08743_ _08744_ _08745_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__nand3_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12863_ _05996_ _05998_ _06029_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__a31oi_2
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _07771_ _07772_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__or2_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _04912_ _05000_ _05001_ _05003_ _04940_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__o221a_1
X_18370_ _02574_ _02588_ _02589_ _02593_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__o31ai_1
XFILLER_15_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _08639_ _08664_ _08669_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__a21o_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _04687_ _04653_ _05645_ _04642_ net34 _05948_ vssd1 vssd1 vccd1 vccd1 _05971_
+ sky130_fd_sc_hd__mux4_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_67_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17321_ _08410_ _08390_ vssd1 vssd1 vccd1 vccd1 _10340_ sky130_fd_sc_hd__and2_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _07686_ _07687_ _07702_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__a21oi_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__buf_4
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _10269_ _10270_ vssd1 vssd1 vccd1 vccd1 _10271_ sky130_fd_sc_hd__nor2_1
XFILLER_187_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14464_ _07634_ _07593_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _04864_ _04865_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a21o_1
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _08373_ _08409_ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__nor2_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13415_ _06585_ _06545_ _06558_ _06564_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__nor4_1
X_10627_ rbzero.tex_r0\[22\] rbzero.tex_r0\[21\] _04099_ vssd1 vssd1 vccd1 vccd1 _04102_
+ sky130_fd_sc_hd__mux2_1
X_17183_ _09542_ _09186_ _10083_ _10202_ vssd1 vssd1 vccd1 vccd1 _10203_ sky130_fd_sc_hd__o31ai_2
X_14395_ _07505_ _07510_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ rbzero.debug_overlay.playerY\[-5\] rbzero.debug_overlay.playerX\[-5\] _08138_
+ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__mux2_1
X_13346_ _06506_ _06488_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__nor2_1
X_10558_ _04065_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16065_ _09155_ _09157_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__and2_1
X_13277_ _06413_ _06436_ _06445_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__and4b_2
X_10489_ _04027_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15016_ net63 _05297_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__nor2_1
X_12228_ rbzero.tex_g1\[27\] _05305_ _05414_ _04947_ vssd1 vssd1 vccd1 vccd1 _05415_
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19824_ rbzero.pov.spi_buffer\[49\] rbzero.pov.spi_buffer\[50\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03524_ sky130_fd_sc_hd__mux2_1
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _04906_ _05344_ _05346_ _04920_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o211a_1
XFILLER_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19670__50 clknet_1_0__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19755_ _03487_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16967_ _09954_ _09988_ vssd1 vssd1 vccd1 vccd1 _09989_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18706_ _02903_ _02904_ _04434_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__o21ai_1
X_15918_ _08253_ _08340_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__or2_1
X_16898_ _09918_ _09919_ vssd1 vssd1 vccd1 vccd1 _09920_ sky130_fd_sc_hd__and2b_1
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ _08335_ _08473_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__nor2_1
X_18637_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__or2_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18568_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__nand2_1
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17519_ _01700_ _01809_ _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a21oi_2
X_18499_ rbzero.map_rom.i_row\[4\] _02718_ _02704_ vssd1 vssd1 vccd1 vccd1 _02719_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22062_ clknet_leaf_79_i_clk _01651_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21013_ clknet_leaf_77_i_clk _00602_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21915_ net441 _01504_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21846_ net372 _01435_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21777_ net303 _01366_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20258__127 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__inv_2
X_11530_ rbzero.map_overlay.i_mapdx\[4\] vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__inv_2
X_20728_ _03934_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__buf_1
XFILLER_157_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20659_ _03734_ _03879_ _03881_ _03740_ rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1
+ _01613_ sky130_fd_sc_hd__a32o_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__mux2_1
X_10412_ rbzero.tex_r1\[57\] rbzero.tex_r1\[58\] _03980_ vssd1 vssd1 vccd1 vccd1 _03987_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14180_ _06854_ _07331_ _07350_ _07336_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__a22oi_2
X_11392_ _04449_ _04581_ _04525_ _04583_ _03971_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a311oi_2
XFILLER_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13131_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__nand2_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ rbzero.map_overlay.i_otherx\[2\] _06120_ rbzero.map_rom.i_row\[4\] _04713_
+ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a22o_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12013_ rbzero.tex_r1\[2\] _05032_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__or2_1
XFILLER_133_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17870_ _02028_ _02065_ _02063_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09848_ sky130_fd_sc_hd__nand2_1
XFILLER_4_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19540_ _03398_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16752_ _09787_ _09788_ vssd1 vssd1 vccd1 vccd1 _09789_ sky130_fd_sc_hd__xnor2_1
X_13964_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__inv_2
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15703_ _08741_ _08785_ _08795_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__a21o_1
X_12915_ _06088_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__and2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16683_ _09749_ vssd1 vssd1 vccd1 vccd1 _09753_ sky130_fd_sc_hd__buf_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19471_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__clkbuf_4
X_13895_ _06718_ _06857_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__nor2_1
X_15634_ _08670_ _08677_ _08676_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__a21o_1
X_18422_ _02635_ _02641_ _02650_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12846_ _06003_ _06021_ _06006_ _06002_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a211o_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _05111_ rbzero.debug_overlay.vplaneX\[-9\] _02576_ vssd1 vssd1 vccd1 vccd1
+ _02587_ sky130_fd_sc_hd__a21oi_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15565_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__or2_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ net44 _05945_ _05941_ net43 _05940_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a221o_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _10189_ _10190_ vssd1 vssd1 vccd1 vccd1 _10323_ sky130_fd_sc_hd__nand2_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _07660_ _07659_ _07651_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__a21o_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19707__84 clknet_1_1__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
X_11728_ _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__buf_6
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18284_ _04432_ _09743_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__or2_1
X_15496_ _08584_ _08589_ _08590_ vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__a21o_1
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _10248_ vssd1 vssd1 vccd1 vccd1 _10255_ sky130_fd_sc_hd__inv_2
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _07603_ _07616_ _07617_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11659_ _04839_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nand2_1
XFILLER_156_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17166_ _10059_ _08553_ _10185_ vssd1 vssd1 vccd1 vccd1 _10186_ sky130_fd_sc_hd__or3_1
XFILLER_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14378_ _07446_ _07478_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__or2_1
XFILLER_196_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16117_ _09165_ _09210_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13329_ _06373_ _06415_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__nand2_1
X_17097_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10118_ sky130_fd_sc_hd__nor2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _09140_ _09141_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__nor2_1
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19807_ rbzero.pov.spi_buffer\[41\] rbzero.pov.spi_buffer\[42\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20363__222 clknet_1_0__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__inv_2
X_17999_ _02137_ _02228_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__nand2_1
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19738_ _03478_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21700_ net226 _01289_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21631_ clknet_leaf_80_i_clk _01220_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
X_21562_ clknet_leaf_90_i_clk _01151_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21493_ net211 _01082_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22045_ clknet_leaf_55_i_clk _01634_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _04277_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12700_ _05830_ _05877_ _05878_ _05298_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__o22a_2
X_13680_ _06840_ _06842_ _06845_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ _04241_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ gpout2.clk_div\[1\] _05808_ _05809_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_
+ sky130_fd_sc_hd__a211o_2
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21829_ net355 _01418_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
X_20562__22 clknet_1_1__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15350_ _08144_ _08442_ _08444_ vssd1 vssd1 vccd1 vccd1 _08445_ sky130_fd_sc_hd__o21ai_4
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12562_ _05702_ _05740_ _05742_ net13 vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__o211a_1
XFILLER_145_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14301_ _07467_ _07469_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__xor2_1
XFILLER_141_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11513_ _04683_ _04690_ _04694_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a31o_1
XFILLER_196_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15281_ _08372_ _08374_ _08375_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12493_ _05053_ _05638_ _05663_ _05673_ _05674_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a311o_1
XFILLER_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17020_ _09146_ _09252_ _09915_ _09914_ vssd1 vssd1 vccd1 vccd1 _10041_ sky130_fd_sc_hd__o31ai_2
XFILLER_184_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14232_ _07397_ _07400_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__nand2_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _07067_ _06759_ _07331_ _07307_ _07329_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__a311o_1
X_11375_ _04555_ _04566_ _04449_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__mux2_1
XFILLER_180_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13114_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
XFILLER_125_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18971_ rbzero.spi_registers.spi_buffer\[16\] rbzero.spi_registers.spi_buffer\[15\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__mux2_1
X_14094_ _07220_ _07261_ _07263_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nand3_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _02186_ _02116_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__o21a_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _06120_ _06086_ rbzero.map_rom.a6 _06219_ _06220_ vssd1 vssd1 vccd1 vccd1
+ _06221_ sky130_fd_sc_hd__a2111o_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17853_ _02140_ _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__xor2_1
XFILLER_94_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16804_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09833_ sky130_fd_sc_hd__nand2_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17784_ _02070_ _02072_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__and2_1
X_14996_ rbzero.wall_tracer.stepDistX\[3\] _08006_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08108_ sky130_fd_sc_hd__mux2_1
XFILLER_94_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19523_ _03389_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13947_ _06942_ _06718_ _07116_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__o21ai_1
X_16735_ rbzero.map_rom.f1 _09118_ vssd1 vssd1 vccd1 vccd1 _09773_ sky130_fd_sc_hd__or2_1
XFILLER_35_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19454_ rbzero.spi_registers.new_vshift\[1\] _02481_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03353_ sky130_fd_sc_hd__mux2_1
X_16666_ _09744_ vssd1 vssd1 vccd1 vccd1 _09745_ sky130_fd_sc_hd__clkbuf_4
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _07034_ _07035_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__nand2_1
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ _08213_ _08250_ _08251_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__or3b_1
X_18405_ _02597_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02635_
+ sky130_fd_sc_hd__nand2_1
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _06003_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__and2_1
X_16597_ _06433_ _08338_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__nor2_2
X_19385_ _03313_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ _08642_ _08236_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__xnor2_1
X_18336_ _02569_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _02571_
+ sky130_fd_sc_hd__and2_1
XFILLER_124_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18267_ _02508_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__clkbuf_1
X_15479_ _08505_ _08506_ _08512_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__a21o_1
XFILLER_129_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _10236_ _10237_ vssd1 vssd1 vccd1 vccd1 _10238_ sky130_fd_sc_hd__nor2_1
XFILLER_129_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18198_ _02462_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__nor2_1
XFILLER_156_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17149_ _10167_ _10165_ vssd1 vssd1 vccd1 vccd1 _10169_ sky130_fd_sc_hd__and2b_1
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03787_ clknet_0__03787_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03787_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20160_ _03728_ _03743_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__and3_1
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20091_ rbzero.pov.ready_buffer\[19\] _03684_ _03699_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01227_ sky130_fd_sc_hd__o211a_1
XFILLER_44_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ clknet_leaf_2_i_clk _00582_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21614_ clknet_leaf_89_i_clk _01203_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_205_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21545_ clknet_leaf_71_i_clk _01134_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21476_ net194 _01065_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11160_ _04381_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11091_ _04345_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22028_ clknet_leaf_55_i_clk _01617_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ rbzero.wall_tracer.stepDistY\[3\] _08006_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08007_ sky130_fd_sc_hd__mux2_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _06966_ _06968_ _06967_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__o21ai_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14781_ _06577_ _07855_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__or2_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11993_ _04830_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__buf_4
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16520_ _09607_ _09609_ vssd1 vssd1 vccd1 vccd1 _09610_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13732_ _06729_ _06758_ _06901_ _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nand4_2
X_10944_ _04268_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20500__346 clknet_1_0__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__inv_2
XFILLER_188_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _09406_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__clkbuf_4
X_13663_ _06832_ _06833_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__xor2_1
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10875_ _04232_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _08400_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _05711_ _05793_ net50 vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a21oi_1
X_19170_ _03175_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__buf_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _09472_ _09473_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13594_ _06762_ _06763_ _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__and3_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _02394_ _02395_ _02396_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a21oi_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _08424_ _08427_ _08161_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__a21o_2
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ net13 _05703_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nor2_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18052_ _09872_ _02334_ _02335_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__o31a_1
XFILLER_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15264_ _08340_ _08358_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__or2_1
XFILLER_177_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12476_ net4 vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__inv_2
XFILLER_172_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17003_ _09929_ _09994_ vssd1 vssd1 vccd1 vccd1 _10024_ sky130_fd_sc_hd__nand2_1
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14215_ _07345_ _07346_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
XANTENNA_5 _05064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ rbzero.spi_registers.texadd0\[0\] _04535_ _04618_ _03970_ vssd1 vssd1 vccd1
+ vccd1 _04619_ sky130_fd_sc_hd__o211a_1
X_15195_ _08238_ _08289_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _07305_ _07315_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__xor2_1
XFILLER_126_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ rbzero.spi_registers.texadd3\[21\] _04526_ _04537_ rbzero.spi_registers.texadd2\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a22o_1
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14077_ _07212_ _07247_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__xnor2_4
X_18954_ rbzero.spi_registers.spi_buffer\[8\] rbzero.spi_registers.spi_buffer\[7\]
+ _03052_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11289_ rbzero.texu_hot\[4\] _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__nand2_1
X_17905_ _02191_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__xnor2_1
X_13028_ _06178_ _06203_ _06176_ _06177_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18885_ rbzero.pov.spi_buffer\[50\] rbzero.pov.ready_buffer\[50\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _10315_ _09363_ _02124_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or3_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ _02054_ _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__xor2_1
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14979_ rbzero.wall_tracer.stepDistX\[-5\] _07954_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08099_ sky130_fd_sc_hd__mux2_1
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19506_ _03379_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__clkbuf_4
X_16718_ _09751_ vssd1 vssd1 vccd1 vccd1 _09759_ sky130_fd_sc_hd__buf_2
X_17698_ _01986_ _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nor2_1
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19437_ _03343_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
X_16649_ _04446_ _04448_ _09735_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a21oi_1
X_20475__323 clknet_1_1__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__inv_2
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ rbzero.spi_registers.new_vshift\[3\] _03297_ _03303_ _03302_ vssd1 vssd1
+ vccd1 vccd1 _00900_ sky130_fd_sc_hd__o211a_1
XFILLER_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _02534_ _02554_ _02555_ _09745_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a31o_1
XFILLER_187_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19299_ rbzero.spi_registers.texadd3\[17\] _03255_ vssd1 vssd1 vccd1 vccd1 _03263_
+ sky130_fd_sc_hd__or2_1
XFILLER_148_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21330_ clknet_leaf_33_i_clk _00919_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21261_ clknet_leaf_3_i_clk _00850_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20212_ rbzero.spi_registers.new_texadd\[3\]\[21\] rbzero.spi_registers.spi_buffer\[21\]
+ _03384_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__mux2_1
X_21192_ clknet_leaf_21_i_clk _00781_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20143_ _09729_ _03092_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__a21bo_1
XFILLER_132_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20074_ rbzero.debug_overlay.vplaneX\[-9\] _03676_ _03690_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01219_ sky130_fd_sc_hd__a211o_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20976_ clknet_leaf_63_i_clk _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ rbzero.tex_r0\[6\] rbzero.tex_r0\[5\] _04110_ vssd1 vssd1 vccd1 vccd1 _04119_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _04077_ vssd1 vssd1 vccd1 vccd1 _04083_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12330_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04908_ vssd1 vssd1 vccd1 vccd1 _05516_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21528_ clknet_leaf_97_i_clk _01117_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ rbzero.tex_g1\[37\] _04817_ _04830_ _04814_ vssd1 vssd1 vccd1 vccd1 _05448_
+ sky130_fd_sc_hd__a31o_1
X_21459_ net177 _01048_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14000_ _06723_ _06738_ _06993_ _06718_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a211o_1
X_11212_ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__clkbuf_8
X_12192_ _05300_ _05378_ _05379_ _04661_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a31o_1
XFILLER_150_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ _04372_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__buf_2
XFILLER_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11074_ _04336_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
X_15951_ rbzero.wall_tracer.stepDistX\[3\] _09045_ vssd1 vssd1 vccd1 vccd1 _09046_
+ sky130_fd_sc_hd__nand2_8
XFILLER_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14902_ rbzero.wall_tracer.visualWallDist\[-9\] _08047_ vssd1 vssd1 vccd1 vccd1 _08048_
+ sky130_fd_sc_hd__or2_1
X_15882_ _08932_ _08934_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__or2_1
X_18670_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__or2_1
XFILLER_62_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__and2_1
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14833_ rbzero.wall_tracer.stepDistY\[0\] _07992_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _07993_ sky130_fd_sc_hd__mux2_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20424__277 clknet_1_1__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__inv_2
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _01726_ _01733_ _01731_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a21oi_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _07067_ _07855_ _06663_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__a21o_1
XFILLER_189_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ rbzero.debug_overlay.playerY\[-6\] _05121_ _05117_ rbzero.debug_overlay.playerY\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a22o_1
XFILLER_189_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13715_ _06876_ _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__xnor2_1
X_16503_ rbzero.debug_overlay.playerY\[-2\] rbzero.debug_overlay.playerX\[-2\] _08138_
+ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__mux2_1
X_10927_ rbzero.tex_g0\[8\] rbzero.tex_g0\[7\] _04259_ vssd1 vssd1 vccd1 vccd1 _04260_
+ sky130_fd_sc_hd__mux2_1
X_17483_ _09647_ _09243_ _09363_ _09519_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__o22a_1
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14695_ _06379_ _06505_ _06515_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__a21o_4
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19222_ rbzero.spi_registers.texadd2\[8\] _03208_ vssd1 vssd1 vccd1 vccd1 _03219_
+ sky130_fd_sc_hd__or2_1
X_16434_ _08731_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__buf_2
XFILLER_147_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13646_ _06763_ _06764_ _06762_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__a21oi_1
X_10858_ _04223_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _09384_ _09456_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ rbzero.spi_registers.new_texadd\[1\]\[2\] _03174_ _03179_ _03169_ vssd1 vssd1
+ vccd1 vccd1 _00809_ sky130_fd_sc_hd__o211a_1
X_13577_ _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__clkbuf_4
X_10789_ rbzero.tex_g1\[8\] rbzero.tex_g1\[9\] _04177_ vssd1 vssd1 vccd1 vccd1 _04187_
+ sky130_fd_sc_hd__mux2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15316_ _08390_ _08400_ _08409_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__o22a_1
X_18104_ _02380_ _02381_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a21oi_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12528_ net14 _05705_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a21oi_1
X_16296_ _08151_ _08165_ _08734_ _08731_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__or4_1
XFILLER_173_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19084_ rbzero.spi_registers.new_mapd\[0\] _03119_ _03138_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00781_ sky130_fd_sc_hd__o211a_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20318__182 clknet_1_1__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__inv_2
XFILLER_184_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15247_ _08331_ _08341_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__xnor2_1
X_18035_ _02245_ _02250_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__or2b_1
X_12459_ net5 _05640_ net7 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a21o_1
XFILLER_160_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ _08160_ _08272_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__nor2_1
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ _07299_ _07255_ _07283_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__o21a_1
XFILLER_98_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19986_ rbzero.debug_overlay.playerY\[-1\] _03611_ _03631_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01190_ sky130_fd_sc_hd__a211o_1
XFILLER_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18937_ _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__buf_4
XFILLER_67_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18868_ rbzero.pov.spi_buffer\[42\] rbzero.pov.ready_buffer\[42\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03015_ sky130_fd_sc_hd__mux2_1
X_17819_ _02106_ _02107_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18799_ rbzero.pov.spi_buffer\[9\] rbzero.pov.ready_buffer\[9\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02979_ sky130_fd_sc_hd__mux2_1
X_20830_ clknet_leaf_50_i_clk _00419_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20761_ _02519_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20692_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03909_
+ sky130_fd_sc_hd__nand2_1
XFILLER_189_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21313_ clknet_leaf_35_i_clk _00902_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21244_ clknet_leaf_26_i_clk _00833_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21175_ clknet_leaf_14_i_clk _00764_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20126_ _04731_ _03719_ _05648_ _03091_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__or4b_1
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20057_ rbzero.debug_overlay.facingY\[-4\] _03658_ vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__or2_1
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ rbzero.row_render.wall\[0\] rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1
+ vccd1 _05020_ sky130_fd_sc_hd__or2b_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04934_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20959_ clknet_leaf_64_i_clk _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _06662_ _06667_ _06670_ _06611_ _06525_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a32o_1
XFILLER_187_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10712_ rbzero.tex_g1\[45\] rbzero.tex_g1\[46\] _04144_ vssd1 vssd1 vccd1 vccd1 _04147_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14480_ _07632_ _07650_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__xnor2_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _03976_ _04864_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__or2_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _06537_ _06539_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__nand2_4
X_10643_ _04054_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16150_ _09242_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__buf_4
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13362_ _06506_ _06488_ _06436_ _06445_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__and4bb_1
X_10574_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _04066_ vssd1 vssd1 vccd1 vccd1 _04074_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15101_ _07866_ _07958_ _07963_ _08143_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__a31o_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ _05497_ _05498_ _04891_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__mux2_1
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ _09166_ _09174_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__xnor2_2
XFILLER_158_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ _06414_ _06417_ _06450_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a21o_1
XFILLER_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _08124_ _08033_ rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__a21o_1
X_12244_ rbzero.tex_g1\[60\] _04904_ _04964_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19840_ rbzero.pov.spi_buffer\[57\] rbzero.pov.spi_buffer\[58\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
X_12175_ _05361_ _05362_ _04947_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__mux2_1
XFILLER_123_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11126_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _04362_ vssd1 vssd1 vccd1 vccd1 _04364_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19771_ rbzero.pov.spi_buffer\[24\] rbzero.pov.spi_buffer\[25\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
X_16983_ _10003_ _10004_ vssd1 vssd1 vccd1 vccd1 _10005_ sky130_fd_sc_hd__and2_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18722_ _02889_ _02907_ _02911_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a21oi_1
X_15934_ _08385_ _09027_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__a21bo_1
X_11057_ rbzero.tex_b1\[9\] rbzero.tex_b1\[10\] _04325_ vssd1 vssd1 vccd1 vccd1 _04328_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _02854_ _02855_ _02841_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a21oi_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _08921_ _08925_ vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17604_ _01700_ _01809_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nand2_1
X_14816_ _07822_ _07807_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__or2_1
XFILLER_188_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18584_ rbzero.debug_overlay.vplaneY\[-5\] _02791_ vssd1 vssd1 vccd1 vccd1 _02792_
+ sky130_fd_sc_hd__xor2_1
Xtop_ew_algofoogle_110 vssd1 vssd1 vccd1 vccd1 ones[1] top_ew_algofoogle_110/LO sky130_fd_sc_hd__conb_1
X_15796_ _08838_ _08890_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__or2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_121 vssd1 vssd1 vccd1 vccd1 ones[12] top_ew_algofoogle_121/LO sky130_fd_sc_hd__conb_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17535_ _01808_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__xor2_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11959_ _05146_ _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__or2_1
X_14747_ _07885_ _07882_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__nor2_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17466_ _01754_ _01756_ _01758_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__o21ai_4
X_14678_ _07842_ _07834_ _07846_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19205_ rbzero.spi_registers.new_texadd\[2\]\[0\] _03206_ _03209_ _03197_ vssd1 vssd1
+ vccd1 vccd1 _00831_ sky130_fd_sc_hd__o211a_1
X_16417_ _09376_ _09496_ _09506_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__and3_1
X_13629_ _06742_ _06743_ _06733_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17397_ _10387_ _01663_ _01688_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__nand3_1
XFILLER_73_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19136_ _03110_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__clkbuf_4
X_16348_ _09313_ _09317_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__and2_1
XFILLER_145_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16279_ _08274_ _08617_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__nor2_1
X_19067_ _03110_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__buf_2
XFILLER_160_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18018_ _10315_ _09890_ _01898_ _09315_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a211oi_1
XFILLER_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19969_ _08223_ rbzero.pov.ready_buffer\[47\] _03561_ vssd1 vssd1 vccd1 vccd1 _03620_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21931_ net457 _01520_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21862_ net388 _01451_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20813_ clknet_leaf_58_i_clk _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21793_ net319 _01382_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20744_ rbzero.traced_texVinit\[9\] _02606_ _03937_ _10126_ vssd1 vssd1 vccd1 vccd1
+ _01643_ sky130_fd_sc_hd__a22o_1
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20675_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03895_
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19656__37 clknet_1_0__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21227_ clknet_leaf_24_i_clk _00816_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21158_ clknet_leaf_12_i_clk _00747_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20109_ rbzero.debug_overlay.vplaneY\[-3\] _03685_ vssd1 vssd1 vccd1 vccd1 _03709_
+ sky130_fd_sc_hd__or2_1
XFILLER_59_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13980_ _07104_ _06888_ _06927_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__or3_1
X_21089_ clknet_leaf_97_i_clk _00678_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12931_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__inv_2
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15650_ _08678_ _08729_ _08742_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__a21o_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12862_ _06031_ _06030_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__and2b_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ rbzero.tex_r0\[50\] _05002_ _04934_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a21o_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _07727_ _07750_ _07749_ _07751_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a22oi_1
XFILLER_2_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15581_ _08671_ _08675_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__xnor2_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _04731_ _05958_ _05948_ _05969_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a211o_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _10329_ _10338_ vssd1 vssd1 vccd1 vccd1 _10339_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14532_ _07686_ _07687_ _07702_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__and3_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11744_ _04891_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__buf_4
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17251_ _10266_ _10267_ _10268_ vssd1 vssd1 vccd1 vccd1 _10270_ sky130_fd_sc_hd__and3_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14463_ _07316_ _07158_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__or2_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11675_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] rbzero.row_render.size\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nand3_1
X_20536__378 clknet_1_1__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__inv_2
X_16202_ _09170_ _09293_ _09294_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__a21o_1
XFILLER_169_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13414_ _06510_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__inv_2
X_10626_ _04101_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__clkbuf_1
X_17182_ _10077_ _10082_ vssd1 vssd1 vccd1 vccd1 _10202_ sky130_fd_sc_hd__nand2_1
X_14394_ _07558_ _07563_ _07564_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__a21bo_1
XFILLER_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16133_ _09125_ _09226_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__xnor2_4
X_13345_ _06379_ _06505_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a21oi_4
X_10557_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _04055_ vssd1 vssd1 vccd1 vccd1 _04065_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16064_ _09155_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__nor2_1
XFILLER_115_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13276_ _06423_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__xor2_1
X_10488_ rbzero.tex_r1\[21\] rbzero.tex_r1\[22\] _04024_ vssd1 vssd1 vccd1 vccd1 _04027_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15015_ _08118_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
X_12227_ rbzero.tex_g1\[26\] _04831_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or2_1
XFILLER_170_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19823_ _03467_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__clkbuf_4
X_12158_ _04923_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__or2_1
XFILLER_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11109_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _04351_ vssd1 vssd1 vccd1 vccd1 _04355_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ rbzero.pov.spi_buffer\[16\] rbzero.pov.spi_buffer\[17\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03487_ sky130_fd_sc_hd__mux2_1
XFILLER_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16966_ _09985_ _09987_ vssd1 vssd1 vccd1 vccd1 _09988_ sky130_fd_sc_hd__xnor2_1
X_12089_ _04741_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nor2_1
X_18705_ _02887_ _02894_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__and2b_1
X_15917_ _08557_ _09011_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16897_ _09912_ _09917_ vssd1 vssd1 vccd1 vccd1 _09919_ sky130_fd_sc_hd__or2_1
X_20281__148 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__inv_2
XFILLER_65_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18636_ _02828_ _02826_ _02814_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__o21ai_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _08431_ _08696_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__nor2_1
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18567_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__or2_1
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15779_ _08298_ _08441_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__nor2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17518_ _10288_ _09662_ _09670_ _01697_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__o22a_1
XFILLER_177_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18498_ rbzero.debug_overlay.playerY\[4\] _02717_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02718_ sky130_fd_sc_hd__mux2_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ _01692_ _01741_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19119_ rbzero.spi_registers.texadd0\[12\] _03156_ vssd1 vssd1 vccd1 vccd1 _03160_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22061_ clknet_leaf_76_i_clk _01650_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21012_ clknet_leaf_76_i_clk _00601_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21914_ net440 _01503_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20340__201 clknet_1_1__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__inv_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21845_ net371 _01434_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21776_ net302 _01365_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20727_ _03728_ clknet_1_1__leaf__05879_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__and2_2
XFILLER_141_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11460_ _04641_ _04644_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nor3_4
XFILLER_184_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20658_ _03880_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__inv_2
XFILLER_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10411_ _03986_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11391_ _04473_ _04513_ _04516_ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o31a_1
X_20589_ _03821_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__and2b_1
XFILLER_164_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nand2_1
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ rbzero.map_overlay.i_otherx\[0\] vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__inv_2
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12012_ rbzero.tex_r1\[4\] _05185_ _05195_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09847_ sky130_fd_sc_hd__nor2_1
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16751_ rbzero.wall_tracer.mapX\[6\] _09119_ _09779_ vssd1 vssd1 vccd1 vccd1 _09788_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13963_ _06732_ _06719_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__nor2_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15702_ _08776_ _08777_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__xor2_1
X_19470_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__clkbuf_4
X_12914_ _06089_ _06076_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__xnor2_1
X_13894_ _06865_ _06874_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16682_ rbzero.row_render.size\[7\] _09752_ _09750_ _07982_ vssd1 vssd1 vccd1 vccd1
+ _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18421_ _02597_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _02650_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15633_ _08680_ _08692_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__xnor2_1
X_12845_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nand2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _02571_ _02584_ _02583_ _02582_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__o211ai_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15564_ _08367_ _08658_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__xnor2_2
X_12776_ _05946_ net34 _05053_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__and3_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _10320_ _10321_ vssd1 vssd1 vccd1 vccd1 _10322_ sky130_fd_sc_hd__xnor2_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _04790_ _04806_ _04813_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__nor3_4
X_14515_ _07660_ _07651_ _07659_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__nand3_1
X_15495_ _08575_ _08576_ _08583_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__and3_1
X_18283_ rbzero.debug_overlay.vplaneX\[-9\] _02522_ _04433_ vssd1 vssd1 vccd1 vccd1
+ _02523_ sky130_fd_sc_hd__mux2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ _10248_ _10253_ vssd1 vssd1 vccd1 vccd1 _10254_ sky130_fd_sc_hd__nand2_1
XFILLER_174_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14446_ _07604_ _07615_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__nor2_1
X_11658_ rbzero.row_render.size\[4\] _04838_ rbzero.row_render.size\[5\] vssd1 vssd1
+ vccd1 vccd1 _04848_ sky130_fd_sc_hd__o21ai_1
XFILLER_168_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ _04092_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__clkbuf_1
X_17165_ rbzero.wall_tracer.visualWallDist\[2\] _08421_ _10183_ _10061_ _10184_ vssd1
+ vssd1 vccd1 vccd1 _10185_ sky130_fd_sc_hd__a41o_1
X_14377_ _07541_ _07547_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__nor2_1
X_11589_ _04774_ _04777_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16116_ _09207_ _09209_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__xor2_1
XFILLER_171_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _06498_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__clkinv_2
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17096_ _09995_ _09996_ _09998_ vssd1 vssd1 vccd1 vccd1 _10117_ sky130_fd_sc_hd__o21a_1
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16047_ _09021_ _09127_ _09139_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__and3_1
X_13259_ _06415_ _06425_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__a21o_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19806_ _03514_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17998_ _02281_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19737_ rbzero.pov.spi_buffer\[8\] rbzero.pov.spi_buffer\[9\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
X_16949_ rbzero.wall_tracer.stepDistY\[10\] _08405_ vssd1 vssd1 vccd1 vccd1 _09971_
+ sky130_fd_sc_hd__nand2_1
XFILLER_38_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18619_ _02809_ _02813_ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19599_ _03428_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__clkbuf_1
X_21630_ clknet_leaf_83_i_clk _01219_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_80_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21561_ clknet_leaf_90_i_clk _01150_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20512_ clknet_1_0__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__buf_1
XFILLER_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21492_ net210 _01081_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19713__88 clknet_1_0__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_101_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22044_ clknet_leaf_41_i_clk _01633_ vssd1 vssd1 vccd1 vccd1 reg_vsync sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_66_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__05700_ clknet_0__05700_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05700_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ rbzero.tex_b1\[55\] rbzero.tex_b1\[56\] _04270_ vssd1 vssd1 vccd1 vccd1 _04277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10891_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _04237_ vssd1 vssd1 vccd1 vccd1 _04241_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ clknet_leaf_40_i_clk _05791_ _05790_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and3_2
X_21828_ net354 _01417_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12561_ net11 _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__or2_1
X_21759_ net285 _01348_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14300_ _07412_ _07470_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__xor2_1
X_11512_ _04696_ _04697_ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or3_2
X_15280_ _08368_ _08246_ _08371_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__or3_1
XFILLER_157_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ net44 _05664_ _05638_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__and3_1
XFILLER_141_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _07335_ _07340_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__nand3b_2
X_11443_ clknet_leaf_35_i_clk vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_19_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _07328_ _07330_ _07332_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__a21bo_1
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11374_ _04559_ _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__and2_1
XFILLER_166_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18970_ _03069_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__clkbuf_1
X_14093_ _07220_ _07261_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__a21o_1
XFILLER_124_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _02205_ _02206_ _02207_ _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__o2bb2a_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _06113_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20347__207 clknet_1_0__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__inv_2
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17852_ _08476_ _02012_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__nor2_1
XFILLER_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16803_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09832_ sky130_fd_sc_hd__nor2_1
XFILLER_94_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17783_ _02070_ _02072_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__nor2_1
XFILLER_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _08107_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19522_ rbzero.spi_registers.new_texadd\[0\]\[3\] _02485_ _03381_ vssd1 vssd1 vccd1
+ vccd1 _03389_ sky130_fd_sc_hd__mux2_1
X_16734_ _09768_ _09771_ _09769_ vssd1 vssd1 vccd1 vccd1 _09772_ sky130_fd_sc_hd__a21o_1
X_13946_ _06942_ _06718_ _07116_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__or3_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _03352_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
X_16665_ _08134_ _09743_ vssd1 vssd1 vccd1 vccd1 _09744_ sky130_fd_sc_hd__nor2_4
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13877_ _06728_ _06983_ _07044_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__o22a_1
X_18404_ _02634_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _08683_ _08684_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__xnor2_1
X_12828_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or2_1
X_19384_ _02485_ rbzero.spi_registers.new_sky\[3\] _03309_ vssd1 vssd1 vccd1 vccd1
+ _03313_ sky130_fd_sc_hd__mux2_1
X_16596_ _09685_ _09566_ _08458_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__a21oi_2
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18335_ _02569_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _02570_
+ sky130_fd_sc_hd__nor2_1
X_15547_ _08237_ _08214_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__nand2_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _05911_ _05921_ _05909_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__nand3_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20393__249 clknet_1_1__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__inv_2
XFILLER_72_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18266_ rbzero.spi_registers.new_texadd\[2\]\[22\] rbzero.spi_registers.spi_buffer\[22\]
+ _02478_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
X_15478_ _08515_ _08525_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__xnor2_1
X_17217_ _10234_ _10235_ vssd1 vssd1 vccd1 vccd1 _10237_ sky130_fd_sc_hd__and2_1
XFILLER_163_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14429_ _07588_ _07595_ _07597_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__and3_1
X_18197_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__nor2_1
X_17148_ _10165_ _10167_ vssd1 vssd1 vccd1 vccd1 _10168_ sky130_fd_sc_hd__and2b_1
XFILLER_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03786_ clknet_0__03786_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03786_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17079_ _10097_ _10099_ vssd1 vssd1 vccd1 vccd1 _10100_ sky130_fd_sc_hd__xor2_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20090_ rbzero.debug_overlay.vplaneX\[-1\] _03685_ vssd1 vssd1 vccd1 vccd1 _03699_
+ sky130_fd_sc_hd__or2_1
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20287__154 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__inv_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20992_ clknet_leaf_5_i_clk _00581_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21613_ clknet_leaf_89_i_clk _01202_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20452__302 clknet_1_1__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__inv_2
X_21544_ clknet_leaf_71_i_clk _01133_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19698__76 clknet_1_1__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21475_ net193 _01064_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20357_ clknet_1_1__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__buf_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11090_ rbzero.tex_b0\[58\] rbzero.tex_b0\[57\] _04340_ vssd1 vssd1 vccd1 vccd1 _04345_
+ sky130_fd_sc_hd__mux2_1
XFILLER_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22027_ clknet_leaf_55_i_clk _01616_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _06966_ _06969_ _06926_ _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__o211ai_4
XFILLER_112_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11992_ _04910_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__clkbuf_4
X_14780_ _07945_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__clkbuf_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10943_ rbzero.tex_b1\[63\] net51 _04188_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__mux2_1
X_13731_ _06658_ _06738_ _06759_ _06681_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__a22o_1
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16450_ _09515_ _09540_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10874_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _04226_ vssd1 vssd1 vccd1 vccd1 _04232_
+ sky130_fd_sc_hd__mux2_1
X_13662_ _06772_ _06791_ _06786_ _06787_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15401_ _08483_ _08491_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__xnor2_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12613_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nor2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _06740_ _06753_ _06752_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a21o_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16381_ _09347_ _09348_ _09350_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__a21oi_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18120_ _02394_ _02395_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__and3_1
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15332_ _08425_ _08426_ _08144_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__a21o_1
X_12544_ net51 _05719_ _05712_ _05263_ _05717_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a221o_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18051_ _02336_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__buf_4
XFILLER_177_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15263_ rbzero.wall_tracer.stepDistX\[-11\] _08357_ _08171_ vssd1 vssd1 vccd1 vccd1
+ _08358_ sky130_fd_sc_hd__a21boi_2
X_12475_ _05643_ _05647_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17002_ _10021_ _10022_ vssd1 vssd1 vccd1 vccd1 _10023_ sky130_fd_sc_hd__nor2_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14214_ _07383_ _07384_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__nand2_1
X_11426_ rbzero.spi_registers.texadd1\[0\] _04545_ _04536_ _04617_ vssd1 vssd1 vccd1
+ vccd1 _04618_ sky130_fd_sc_hd__a211o_1
X_15194_ _08268_ _08288_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__xnor2_1
XANTENNA_6 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14145_ _07078_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__buf_2
X_11357_ _04544_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nand2_1
XFILLER_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ _07213_ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__xor2_4
X_18953_ _03060_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11288_ rbzero.spi_registers.texadd0\[10\] _04467_ _04478_ _04479_ vssd1 vssd1 vccd1
+ vccd1 _04480_ sky130_fd_sc_hd__o22a_1
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17904_ _01922_ _09195_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__or2_1
X_13027_ _06181_ _06198_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nand2_1
XFILLER_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18884_ _03023_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17835_ _08499_ _09243_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__or2_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ _01814_ _01928_ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__o21a_1
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ _08098_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19505_ _08116_ _02936_ _03350_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__and3_1
X_16717_ rbzero.traced_texa\[9\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a22o_1
X_13929_ _07063_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__xnor2_1
X_17697_ _01870_ _01873_ _01871_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__o21a_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19436_ _02487_ rbzero.spi_registers.new_other\[4\] _03338_ vssd1 vssd1 vccd1 vccd1
+ _03343_ sky130_fd_sc_hd__mux2_1
X_16648_ _09734_ _04636_ vssd1 vssd1 vccd1 vccd1 _09735_ sky130_fd_sc_hd__or2_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19367_ rbzero.spi_registers.vshift\[3\] _03298_ vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__or2_1
XFILLER_37_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16579_ _09668_ vssd1 vssd1 vccd1 vccd1 _09669_ sky130_fd_sc_hd__buf_2
XFILLER_210_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18318_ _05120_ _02544_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__or2_1
XFILLER_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19298_ rbzero.spi_registers.new_texadd\[3\]\[16\] _03254_ _03262_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__o211a_1
XFILLER_176_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _02499_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21260_ clknet_leaf_100_i_clk _00849_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20211_ _03772_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21191_ clknet_leaf_18_i_clk _00780_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20142_ _08116_ _03725_ _09731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a21o_1
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20073_ rbzero.pov.ready_buffer\[11\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__and3_1
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20975_ clknet_leaf_61_i_clk _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10590_ _04082_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21527_ clknet_leaf_97_i_clk _01116_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ rbzero.tex_g1\[39\] _05010_ _05446_ _04946_ vssd1 vssd1 vccd1 vccd1 _05447_
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21458_ net176 _01047_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _04052_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__buf_6
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12191_ _05047_ _04683_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nand2_1
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21389_ clknet_leaf_11_i_clk _00978_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _04362_ vssd1 vssd1 vccd1 vccd1 _04372_
+ sky130_fd_sc_hd__mux2_1
XFILLER_134_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__buf_2
XFILLER_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11073_ rbzero.tex_b1\[1\] rbzero.tex_b1\[2\] _03979_ vssd1 vssd1 vccd1 vccd1 _04336_
+ sky130_fd_sc_hd__mux2_1
X_15950_ _08357_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__buf_6
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14901_ _08046_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__buf_2
XFILLER_163_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _08912_ _08943_ _08975_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__and3_1
XFILLER_130_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__nor2_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _06655_ _07988_ _07990_ _07991_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__a211o_4
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _01838_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14763_ _07903_ _07929_ _06669_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__a21oi_1
X_20459__308 clknet_1_1__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__inv_2
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ rbzero.debug_overlay.playerY\[2\] _05103_ _05115_ rbzero.debug_overlay.playerY\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a22o_1
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _09479_ _09592_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__xor2_4
Xclkbuf_1_0__f__03789_ clknet_0__03789_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03789_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ _06779_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17482_ _01714_ _01694_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__or2b_1
X_10926_ _04214_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__buf_4
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14694_ _06568_ _07825_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__o21ba_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ rbzero.spi_registers.new_texadd\[2\]\[7\] _03206_ _03218_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00838_ sky130_fd_sc_hd__o211a_1
X_16433_ _09521_ _09523_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__nand2_1
XFILLER_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10857_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _04215_ vssd1 vssd1 vccd1 vccd1 _04223_
+ sky130_fd_sc_hd__mux2_1
XFILLER_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13645_ _06803_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__and2_1
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ rbzero.spi_registers.texadd1\[2\] _03176_ vssd1 vssd1 vccd1 vccd1 _03179_
+ sky130_fd_sc_hd__or2_1
X_16364_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__nor2_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _04186_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13576_ _06682_ _06693_ _06700_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__and3_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18103_ _02372_ _02375_ _02373_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__o21ai_1
X_15315_ _08213_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_121_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19083_ rbzero.mapdyw\[0\] _03121_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or2_1
X_12527_ _05704_ _05057_ _05706_ net13 _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__o2111a_1
X_16295_ _08151_ _08734_ _08731_ _08166_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__o22ai_1
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _02296_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__xnor2_1
X_15246_ _08337_ _08340_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__or2_1
X_12458_ net6 vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__buf_2
XFILLER_126_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ _04452_ _04584_ _04588_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o31ai_1
X_12389_ _04902_ _05569_ _05573_ _04886_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o31a_1
X_15177_ _04463_ _06063_ _08143_ _08271_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__o211a_1
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14128_ _07257_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__inv_2
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19985_ rbzero.pov.ready_buffer\[52\] _03436_ _03582_ _08322_ _03617_ vssd1 vssd1
+ vccd1 vccd1 _03631_ sky130_fd_sc_hd__o221a_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18936_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__clkbuf_4
X_14059_ _07227_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__and2_1
XFILLER_86_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18867_ _03014_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17818_ _01818_ _10215_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor2_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18798_ _02967_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__clkbuf_4
XFILLER_208_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17749_ _02037_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__nor2_1
XFILLER_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20325__187 clknet_1_1__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__inv_2
XFILLER_208_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20399__255 clknet_1_0__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__inv_2
X_20760_ _05120_ rbzero.wall_tracer.rayAddendX\[-6\] vssd1 vssd1 vccd1 vccd1 _03947_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19419_ _03333_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20691_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03908_
+ sky130_fd_sc_hd__or2_1
XFILLER_210_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21312_ clknet_leaf_34_i_clk _00901_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21243_ clknet_leaf_26_i_clk _00832_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21174_ clknet_leaf_14_i_clk _00763_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20125_ _05651_ _05650_ _05644_ _04687_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or4bb_1
XFILLER_132_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20056_ rbzero.debug_overlay.facingY\[-5\] _03676_ _03679_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01212_ sky130_fd_sc_hd__a211o_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _04908_ vssd1 vssd1 vccd1 vccd1 _04950_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ clknet_leaf_64_i_clk _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _04146_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ rbzero.row_render.size\[9\] _04864_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_
+ sky130_fd_sc_hd__o21a_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ clknet_leaf_46_i_clk _00478_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10642_ _04109_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__clkbuf_1
X_13430_ _06598_ _06599_ _06600_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__a21o_1
XFILLER_167_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _06458_ _06531_ _06518_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__o21ai_1
X_10573_ _04073_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15100_ _08194_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__buf_2
X_12312_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _04907_ vssd1 vssd1 vccd1 vccd1 _05498_
+ sky130_fd_sc_hd__mux2_1
X_16080_ _09169_ _09173_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__xnor2_1
X_13292_ _06332_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__xnor2_4
XFILLER_182_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12243_ rbzero.tex_g1\[61\] _04891_ _04830_ _04814_ vssd1 vssd1 vccd1 vccd1 _05430_
+ sky130_fd_sc_hd__a31o_1
X_15031_ _08128_ rbzero.mapdxw\[0\] _06151_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__mux2_1
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _04964_ vssd1 vssd1 vccd1 vccd1 _05362_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11125_ _04363_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
X_19770_ _03495_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
X_16982_ _09891_ _10002_ vssd1 vssd1 vccd1 vccd1 _10004_ sky130_fd_sc_hd__or2_1
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18721_ _02916_ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__xnor2_1
X_15933_ _08369_ _08408_ _08384_ _08516_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__o22ai_1
X_11056_ _04327_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18652_ _02844_ _02847_ _02853_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__nand3_1
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _08947_ _08957_ _08958_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__or3_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _10059_ _09252_ _01790_ _01788_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__o31ai_2
XFILLER_188_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _07976_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _05129_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.debug_overlay.vplaneY\[-8\]
+ _02756_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__o31a_1
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_100 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_100/HI zeros[7] sky130_fd_sc_hd__conb_1
X_15795_ _08889_ _08344_ _08696_ _08516_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__o22a_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_111 vssd1 vssd1 vccd1 vccd1 ones[2] top_ew_algofoogle_111/LO sky130_fd_sc_hd__conb_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_122 vssd1 vssd1 vccd1 vccd1 ones[13] top_ew_algofoogle_122/LO sky130_fd_sc_hd__conb_1
X_17534_ _01813_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__xnor2_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _07878_ _07884_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__nor2_1
X_11958_ rbzero.debug_overlay.facingX\[-6\] _05121_ _05118_ rbzero.debug_overlay.facingX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a22o_1
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17465_ _01754_ _01756_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a21oi_1
X_10909_ _04250_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ _07847_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__inv_2
X_11889_ _05077_ _05061_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__or2b_1
X_19204_ rbzero.spi_registers.texadd2\[0\] _03208_ vssd1 vssd1 vccd1 vccd1 _03209_
+ sky130_fd_sc_hd__or2_1
X_16416_ _09376_ _09496_ _09506_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _06640_ _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nor2_1
X_17396_ _10387_ _01663_ _01688_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__a21o_1
XFILLER_158_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19135_ rbzero.spi_registers.texadd0\[20\] _03142_ vssd1 vssd1 vccd1 vccd1 _03168_
+ sky130_fd_sc_hd__or2_1
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ _09436_ _09437_ _09420_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__a21o_1
XFILLER_201_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13559_ _06658_ _06729_ _06681_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__a21oi_2
XFILLER_186_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19066_ rbzero.map_overlay.i_mapdy\[0\] _03122_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or2_1
X_16278_ _08296_ _09076_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__nor2_1
X_20513__357 clknet_1_0__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__inv_2
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ _09315_ _01898_ _09890_ _10315_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__o211a_1
XFILLER_173_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ rbzero.wall_tracer.visualWallDist\[-1\] _08158_ _08319_ _08323_ vssd1 vssd1
+ vccd1 vccd1 _08324_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19968_ rbzero.debug_overlay.playerY\[-7\] _03617_ _03619_ _03579_ vssd1 vssd1 vccd1
+ vccd1 _01184_ sky130_fd_sc_hd__o211a_1
XFILLER_68_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18919_ _03041_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19899_ _03559_ _03564_ _03566_ _03302_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__o211a_1
XFILLER_68_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21930_ net456 _01519_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20407__262 clknet_1_0__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__inv_2
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21861_ net387 _01450_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20812_ clknet_leaf_58_i_clk _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21792_ net318 _01381_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20743_ rbzero.traced_texVinit\[8\] _09759_ _03937_ _10010_ vssd1 vssd1 vccd1 vccd1
+ _01642_ sky130_fd_sc_hd__a22o_1
XFILLER_169_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20674_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03894_
+ sky130_fd_sc_hd__nor2_1
XFILLER_195_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21226_ clknet_leaf_24_i_clk _00815_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21157_ clknet_leaf_12_i_clk _00746_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20108_ _05132_ _03655_ _03708_ _03695_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a211o_1
X_21088_ clknet_leaf_97_i_clk _00677_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20039_ rbzero.pov.ready_buffer\[40\] _03656_ _03670_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01204_ sky130_fd_sc_hd__o211a_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _04429_ _04430_ rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__nor3b_2
XFILLER_207_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12861_ _06032_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__xor2_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _07728_ _07730_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04978_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__buf_4
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _08673_ _08674_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__and2_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _05648_ _05958_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nor2_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14531_ _07689_ _07700_ _07701_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a21bo_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__buf_4
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _10266_ _10267_ _10268_ vssd1 vssd1 vccd1 vccd1 _10269_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14462_ _07252_ _07361_ _07632_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__or3_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] rbzero.row_render.size\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a21o_1
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16201_ _08516_ _08400_ _08429_ _08369_ vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__o22a_1
XFILLER_186_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13413_ _06554_ _06578_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__xnor2_4
X_17181_ _10180_ _10200_ vssd1 vssd1 vccd1 vccd1 _10201_ sky130_fd_sc_hd__xor2_1
X_10625_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _04099_ vssd1 vssd1 vccd1 vccd1 _04101_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14393_ _07560_ _07562_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__or2b_1
XFILLER_195_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _09126_ _09225_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__xor2_4
X_10556_ _04064_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13344_ _06507_ _06480_ _06514_ _06467_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__or4b_4
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _08253_ _08535_ _09012_ _09156_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__o31a_1
XFILLER_155_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10487_ _04026_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _06330_ _06431_ _06411_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a21oi_2
XFILLER_182_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ _08117_ _05057_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__and2_1
X_12226_ rbzero.tex_g1\[28\] _04905_ _05305_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _05002_ vssd1 vssd1 vccd1 vccd1 _05345_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19822_ _03522_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _04354_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16965_ _09676_ _09700_ _09986_ vssd1 vssd1 vccd1 vccd1 _09987_ sky130_fd_sc_hd__a21bo_1
X_19753_ _03486_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
X_12088_ _04579_ _05269_ _05271_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__o31a_1
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15916_ _08370_ _08328_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__nor2_1
X_11039_ _04318_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
X_18704_ _02822_ rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 _02903_
+ sky130_fd_sc_hd__xnor2_1
X_16896_ _09912_ _09917_ vssd1 vssd1 vccd1 vccd1 _09918_ sky130_fd_sc_hd__and2_1
XFILLER_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18635_ _02826_ _02829_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__nand2_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _08906_ _08941_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ rbzero.wall_tracer.rayAddendY\[-3\] _02527_ _02772_ _02775_ vssd1 vssd1 vccd1
+ vccd1 _00626_ sky130_fd_sc_hd__o22a_1
X_15778_ _08846_ _08872_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__xor2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17517_ _10288_ _09670_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__nor2_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14729_ _07820_ _07815_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__nand2_1
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18497_ _02716_ _06097_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _01738_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__xor2_1
XFILLER_162_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _01670_ _01671_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__xor2_1
XFILLER_146_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20437__288 clknet_1_0__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__inv_2
XFILLER_158_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19118_ rbzero.spi_registers.new_texadd\[0\]\[11\] _03155_ _03159_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__o211a_1
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20390_ clknet_1_0__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__buf_1
XFILLER_161_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19049_ rbzero.spi_registers.new_vinf _03115_ _03116_ _03117_ _03118_ vssd1 vssd1
+ vccd1 vccd1 _00766_ sky130_fd_sc_hd__o311a_1
XFILLER_160_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22060_ clknet_leaf_76_i_clk _01649_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21011_ clknet_leaf_77_i_clk _00600_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21913_ net439 _01502_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21844_ net370 _01433_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21775_ net301 _01364_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20726_ _03933_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__buf_1
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20657_ _03876_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__and3_1
XFILLER_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10410_ rbzero.tex_r1\[58\] rbzero.tex_r1\[59\] _03980_ vssd1 vssd1 vccd1 vccd1 _03986_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11390_ _04449_ _04517_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__nor2_1
X_20588_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03822_
+ sky130_fd_sc_hd__nand2_1
XFILLER_104_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ _06234_ rbzero.map_rom.i_col\[4\] _06086_ rbzero.map_overlay.i_othery\[2\]
+ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a221o_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12011_ rbzero.tex_r1\[5\] _05199_ _05032_ _04890_ vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21209_ clknet_leaf_11_i_clk _00798_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16750_ rbzero.wall_tracer.mapX\[7\] _09118_ vssd1 vssd1 vccd1 vccd1 _09787_ sky130_fd_sc_hd__xor2_1
XFILLER_24_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13962_ _07090_ _07132_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__nand2_1
XFILLER_115_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _08741_ _08785_ _08795_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12913_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__clkinv_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16681_ _09751_ vssd1 vssd1 vccd1 vccd1 _09752_ sky130_fd_sc_hd__buf_4
XFILLER_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13893_ _06862_ _06864_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__or2b_1
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18420_ _09753_ _02640_ _02641_ _02649_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a31o_1
X_15632_ _08695_ _08705_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__nand2_1
XFILLER_146_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _02582_ _02583_ _02584_ _02571_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a211o_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _08628_ _08657_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__xor2_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ net37 vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__inv_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _09662_ _09046_ _09397_ vssd1 vssd1 vccd1 vccd1 _10321_ sky130_fd_sc_hd__a21oi_2
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14514_ _07682_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__nor2_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _04912_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__or2_1
XFILLER_187_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18282_ _02512_ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15494_ _08587_ _08588_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__and2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ _10009_ _10249_ _10252_ vssd1 vssd1 vccd1 vccd1 _10253_ sky130_fd_sc_hd__o21ai_2
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14445_ _07604_ _07615_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__xor2_1
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11657_ _04840_ _04846_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nor2_1
XFILLER_174_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10608_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _04088_ vssd1 vssd1 vccd1 vccd1 _04092_
+ sky130_fd_sc_hd__mux2_1
X_17164_ _08165_ _08399_ _08499_ _08151_ vssd1 vssd1 vccd1 vccd1 _10184_ sky130_fd_sc_hd__o22a_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14376_ _07491_ _07543_ _07544_ _07546_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11588_ _04774_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nor2_1
XFILLER_183_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _09035_ _09063_ _09208_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ _06496_ _06497_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__xor2_4
X_17095_ _10023_ _10115_ vssd1 vssd1 vccd1 vccd1 _10116_ sky130_fd_sc_hd__xnor2_1
X_10539_ net49 rbzero.tex_r0\[63\] _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__mux2_1
XFILLER_171_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16046_ _09021_ _09127_ _09139_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__a21oi_1
XFILLER_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ _06324_ _06426_ _06428_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__o21ba_1
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12209_ rbzero.tex_g1\[2\] _04831_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__or2_1
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13189_ rbzero.wall_tracer.visualWallDist\[-4\] _06327_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a21o_1
XFILLER_111_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19805_ rbzero.pov.spi_buffer\[40\] rbzero.pov.spi_buffer\[41\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03514_ sky130_fd_sc_hd__mux2_1
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17997_ _02282_ _02283_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16948_ rbzero.wall_tracer.stepDistX\[10\] _09045_ vssd1 vssd1 vccd1 vccd1 _09970_
+ sky130_fd_sc_hd__nand2_2
X_19736_ _03477_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ _09615_ _09900_ vssd1 vssd1 vccd1 vccd1 _09901_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18618_ _02822_ rbzero.wall_tracer.rayAddendY\[2\] vssd1 vssd1 vccd1 vccd1 _02823_
+ sky130_fd_sc_hd__xnor2_1
X_19598_ rbzero.spi_registers.new_texadd\[1\]\[16\] rbzero.spi_registers.spi_buffer\[16\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18549_ _02743_ _02754_ _02744_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21560_ clknet_leaf_90_i_clk _01149_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20519__363 clknet_1_0__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__inv_2
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21491_ net209 _01080_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20370__228 clknet_1_0__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__inv_2
XFILLER_158_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22043_ clknet_leaf_38_i_clk _01632_ vssd1 vssd1 vccd1 vccd1 reg_hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20264__133 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__inv_2
XFILLER_21_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10890_ _04240_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
X_21827_ net353 _01416_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12560_ _04687_ _04653_ _05645_ _04642_ net10 net12 vssd1 vssd1 vccd1 vccd1 _05741_
+ sky130_fd_sc_hd__mux4_1
X_21758_ net284 _01347_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _03972_ _04698_ _04700_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _04701_
+ sky130_fd_sc_hd__o31a_1
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20709_ _04437_ _09729_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__nand2_1
X_12491_ net46 _05659_ _05638_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a31o_1
X_21689_ net215 _01278_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
X_14230_ _07397_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__or2_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11442_ _04415_ _04426_ _04451_ _04580_ _04633_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__a32o_2
XFILLER_165_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14161_ _07316_ _07306_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__or3_1
X_11373_ _04562_ _04563_ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_1
XFILLER_180_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13112_ _06266_ _06282_ _06283_ _06265_ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1
+ vccd1 vccd1 _00390_ sky130_fd_sc_hd__a32o_1
XFILLER_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _07067_ _06758_ _07219_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__a31o_1
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17920_ _01840_ _02093_ _02205_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nor3_1
XFILLER_140_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _06108_ _06130_ rbzero.map_rom.b6 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1
+ _06219_ sky130_fd_sc_hd__a22o_1
XFILLER_105_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17851_ _02138_ _02139_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__nand2_1
XFILLER_61_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16802_ _06186_ _09786_ _09831_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17782_ _01880_ _01961_ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a21oi_1
X_14994_ rbzero.wall_tracer.stepDistX\[2\] _08000_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08107_ sky130_fd_sc_hd__mux2_1
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16733_ _09769_ _09770_ vssd1 vssd1 vccd1 vccd1 _09771_ sky130_fd_sc_hd__nor2_1
X_19521_ _03388_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
X_13945_ _07067_ _07115_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nand2_1
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19452_ rbzero.spi_registers.new_vshift\[0\] _02473_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03352_ sky130_fd_sc_hd__mux2_1
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16664_ rbzero.trace_state\[0\] _05050_ _09729_ vssd1 vssd1 vccd1 vccd1 _09743_ sky130_fd_sc_hd__and3_2
X_13876_ _07026_ _07027_ _07028_ _07046_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__a211o_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15615_ _08708_ _08709_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__xnor2_2
X_18403_ rbzero.wall_tracer.rayAddendX\[4\] _02633_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_62_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12827_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nand2_1
X_19383_ _03312_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
X_16595_ rbzero.wall_tracer.stepDistY\[9\] _08405_ vssd1 vssd1 vccd1 vccd1 _09685_
+ sky130_fd_sc_hd__nand2_1
XFILLER_188_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18334_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__clkbuf_4
X_15546_ _08635_ _08640_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__xor2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12758_ _05898_ _05907_ _05930_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__or4_2
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ rbzero.floor_leak\[5\] _04810_ _04885_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_
+ sky130_fd_sc_hd__a211oi_1
X_18265_ _02507_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__clkbuf_1
X_15477_ _08528_ _08571_ vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12689_ _05866_ _05867_ _05824_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__mux2_1
X_17216_ _10234_ _10235_ vssd1 vssd1 vccd1 vccd1 _10236_ sky130_fd_sc_hd__nor2_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _07554_ _07571_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__xnor2_1
X_18196_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__and2_1
XFILLER_200_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _09647_ _08620_ _10062_ _10166_ vssd1 vssd1 vccd1 vccd1 _10167_ sky130_fd_sc_hd__o31ai_1
X_14359_ _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03785_ clknet_0__03785_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03785_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17078_ _09968_ _09980_ _10098_ vssd1 vssd1 vccd1 vccd1 _10099_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16029_ _08148_ _09122_ _09123_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__or3_2
XFILLER_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19719_ rbzero.pov.mosi rbzero.pov.spi_buffer\[0\] _03468_ vssd1 vssd1 vccd1 vccd1
+ _03469_ sky130_fd_sc_hd__mux2_1
X_20991_ clknet_leaf_24_i_clk _00580_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21612_ clknet_leaf_89_i_clk _01201_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21543_ clknet_leaf_71_i_clk _01132_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21474_ net192 _01063_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22026_ clknet_leaf_39_i_clk _01615_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _05019_ _05030_ _05177_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a31o_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _06772_ _06754_ _06727_ _06755_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__or4_2
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10942_ _04267_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13661_ _06830_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__xor2_1
X_10873_ _04231_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _08419_ _08494_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__xnor2_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ net17 _05763_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nand2_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _09470_ _09471_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__or2_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _06740_ _06752_ _06753_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__nand3_1
XFILLER_185_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _07992_ _07996_ _08393_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__nand3_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ net40 _05720_ _05715_ net41 vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a22o_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ _08139_ _08405_ _04433_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__o21a_2
X_15262_ _08162_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__buf_4
XFILLER_184_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _05640_ _05649_ _05655_ net5 vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__o211a_1
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17001_ _09926_ _10019_ _10020_ vssd1 vssd1 vccd1 vccd1 _10022_ sky130_fd_sc_hd__and3_1
X_14213_ _07377_ _07374_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__xor2_2
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ rbzero.spi_registers.texadd2\[0\] _04537_ _04457_ rbzero.spi_registers.texadd3\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a22o_1
X_15193_ _08276_ _08287_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__nor2_1
XANTENNA_7 _05552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _06738_ _07310_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__nand2_1
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ rbzero.spi_registers.texadd0\[20\] _04535_ _04547_ vssd1 vssd1 vccd1 vccd1
+ _04548_ sky130_fd_sc_hd__o21a_1
XFILLER_67_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14075_ _07214_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__xnor2_4
X_18952_ rbzero.spi_registers.spi_buffer\[7\] rbzero.spi_registers.spi_buffer\[6\]
+ _03052_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ rbzero.spi_registers.texadd3\[10\] _04465_ _04456_ rbzero.spi_registers.texadd2\[10\]
+ _04470_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a221o_1
X_17903_ _02189_ _02190_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__xnor2_1
X_13026_ rbzero.wall_tracer.trackDistX\[1\] vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__inv_2
XFILLER_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18883_ rbzero.pov.spi_buffer\[49\] rbzero.pov.ready_buffer\[49\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17834_ _02059_ _02042_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or2b_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17765_ _01818_ _09677_ _01929_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__or3_1
X_14977_ rbzero.wall_tracer.stepDistX\[-6\] _07944_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08098_ sky130_fd_sc_hd__mux2_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19504_ rbzero.spi_registers.got_new_mapd _03118_ _03316_ _03362_ vssd1 vssd1 vccd1
+ vccd1 _00961_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_50_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16716_ rbzero.traced_texa\[8\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a22o_1
X_13928_ _07086_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__xor2_1
X_17696_ _01984_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__or2b_1
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19435_ _03342_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
X_16647_ _04408_ vssd1 vssd1 vccd1 vccd1 _09734_ sky130_fd_sc_hd__buf_6
X_13859_ _06978_ _07024_ _07028_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__and3_1
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16578_ _09053_ _09306_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__and2_1
X_19366_ rbzero.spi_registers.new_vshift\[2\] _03297_ _03301_ _03302_ vssd1 vssd1
+ vccd1 vccd1 _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15529_ _08622_ _08623_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__or2_1
XFILLER_163_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18317_ _05120_ _02544_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__nand2_1
X_19297_ rbzero.spi_registers.texadd3\[16\] _03255_ vssd1 vssd1 vccd1 vccd1 _03262_
+ sky130_fd_sc_hd__or2_1
XFILLER_37_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18248_ rbzero.spi_registers.new_texadd\[2\]\[13\] rbzero.spi_registers.spi_buffer\[13\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XFILLER_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__nor2_1
XFILLER_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20210_ rbzero.spi_registers.new_texadd\[3\]\[20\] rbzero.spi_registers.spi_buffer\[20\]
+ _03384_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__mux2_1
X_21190_ clknet_leaf_20_i_clk _00779_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20141_ _03731_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03799_ _03799_ vssd1 vssd1 vccd1 vccd1 clknet_0__03799_ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20072_ rbzero.debug_overlay.facingY\[10\] _03676_ _03689_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01218_ sky130_fd_sc_hd__a211o_1
X_20482__329 clknet_1_0__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__inv_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_18_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ clknet_leaf_61_i_clk _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20376__234 clknet_1_1__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__inv_2
XFILLER_194_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21526_ clknet_leaf_97_i_clk _01115_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21457_ net175 _01046_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
X_11210_ _04407_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__clkbuf_1
X_12190_ _05370_ _05376_ _05377_ _04900_ _04702_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__o221ai_2
X_21388_ clknet_leaf_2_i_clk _00977_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _04371_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__buf_2
X_11072_ _04335_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14900_ _08045_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__buf_2
XFILLER_114_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22009_ clknet_leaf_37_i_clk _01598_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _08973_ _08974_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__xor2_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _06602_ _06598_ _07917_ _06516_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__a31o_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _01841_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__buf_2
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14762_ _07904_ _07901_ _07894_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__mux2_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ rbzero.debug_overlay.playerX\[2\] _05103_ _05155_ _05162_ vssd1 vssd1 vccd1
+ vccd1 _05163_ sky130_fd_sc_hd__a211oi_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _09590_ _09591_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__nand2_2
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03788_ clknet_0__03788_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03788_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13713_ _06882_ _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10925_ _04258_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17481_ _01713_ _01696_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__or2b_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14693_ _07826_ _07862_ _07863_ _06568_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__o211a_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16432_ _08152_ _09520_ _09522_ vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__or3_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19220_ rbzero.spi_registers.texadd2\[7\] _03208_ vssd1 vssd1 vccd1 vccd1 _03218_
+ sky130_fd_sc_hd__or2_1
X_13644_ _06812_ _06813_ _06814_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__a21bo_1
X_10856_ _04222_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ rbzero.spi_registers.new_texadd\[1\]\[1\] _03174_ _03178_ _03169_ vssd1 vssd1
+ vccd1 vccd1 _00808_ sky130_fd_sc_hd__o211a_1
X_16363_ _09452_ _09453_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__and2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13575_ _06745_ _06744_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__xnor2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ rbzero.tex_g1\[9\] rbzero.tex_g1\[10\] _04177_ vssd1 vssd1 vccd1 vccd1 _04186_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__nand2_1
X_15314_ _08408_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__clkbuf_4
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ rbzero.spi_registers.new_mapd\[3\] _03119_ _03137_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00780_ sky130_fd_sc_hd__o211a_1
X_12526_ net14 vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__inv_2
XFILLER_185_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ _09289_ _09299_ _09298_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__a21bo_1
XFILLER_9_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18033_ _02297_ _02319_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _06263_ _08218_ _08315_ _08339_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__o31a_4
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12457_ _05637_ _05638_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nand2_1
XFILLER_138_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11408_ _04589_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__nor2_1
X_15176_ _04463_ _06382_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__nand2_1
XFILLER_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12388_ _05190_ _05570_ _05571_ _05572_ _04940_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__o221a_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14127_ _07242_ _07282_ _07296_ _07280_ _07297_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__a221o_1
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11339_ rbzero.spi_registers.texadd3\[17\] _04526_ _04456_ rbzero.spi_registers.texadd2\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__a22o_1
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19984_ rbzero.debug_overlay.playerY\[-2\] _03617_ _03629_ _03630_ vssd1 vssd1 vccd1
+ vccd1 _01189_ sky130_fd_sc_hd__o211a_1
XFILLER_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18935_ _03049_ _02929_ _02951_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__and3b_1
X_14058_ _07135_ _07225_ _07226_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__o22ai_1
XFILLER_80_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13009_ rbzero.wall_tracer.trackDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__inv_2
XFILLER_140_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18866_ rbzero.pov.spi_buffer\[41\] rbzero.pov.ready_buffer\[41\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17817_ _02050_ _02105_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__xnor2_1
X_18797_ _02977_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17748_ _01842_ _01949_ _01839_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a21boi_1
XFILLER_130_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17679_ _01968_ _01969_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__nand2_1
XFILLER_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19418_ _02485_ rbzero.spi_registers.new_leak\[3\] _03329_ vssd1 vssd1 vccd1 vccd1
+ _03333_ sky130_fd_sc_hd__mux2_1
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20690_ rbzero.texV\[7\] _03814_ _03819_ _03907_ vssd1 vssd1 vccd1 vccd1 _01618_
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19349_ rbzero.color_floor\[1\] _03289_ _03292_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__a21o_1
XFILLER_206_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21311_ clknet_leaf_34_i_clk _00900_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21242_ clknet_leaf_26_i_clk _00831_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21173_ clknet_leaf_22_i_clk _00762_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20124_ _05644_ _03716_ _04691_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__and4_1
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20055_ rbzero.pov.ready_buffer\[26\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__and3_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ clknet_leaf_64_i_clk _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10710_ rbzero.tex_g1\[46\] rbzero.tex_g1\[47\] _04144_ vssd1 vssd1 vccd1 vccd1 _04146_
+ sky130_fd_sc_hd__mux2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ rbzero.row_render.size\[9\] _04864_ _03976_ vssd1 vssd1 vccd1 vccd1 _04880_
+ sky130_fd_sc_hd__a21o_1
XFILLER_201_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20888_ clknet_leaf_44_i_clk _00477_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_1
X_10641_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _04099_ vssd1 vssd1 vccd1 vccd1 _04109_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ _06528_ _06455_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__and2_1
X_10572_ rbzero.tex_r0\[48\] rbzero.tex_r0\[47\] _04066_ vssd1 vssd1 vccd1 vccd1 _04073_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12311_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _04893_ vssd1 vssd1 vccd1 vccd1 _05497_
+ sky130_fd_sc_hd__mux2_1
X_21509_ clknet_leaf_81_i_clk _01098_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _06345_ _06409_ _06411_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a21oi_2
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ rbzero.mapdyw\[0\] _06159_ _08127_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__a21bo_1
XFILLER_170_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12242_ rbzero.tex_g1\[63\] _05010_ _05428_ _04946_ vssd1 vssd1 vccd1 vccd1 _05429_
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _04932_ vssd1 vssd1 vccd1 vccd1 _05361_
+ sky130_fd_sc_hd__mux2_1
X_20430__283 clknet_1_1__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__inv_2
XFILLER_64_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19682__61 clknet_1_1__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
X_11124_ rbzero.tex_b0\[42\] rbzero.tex_b0\[41\] _04362_ vssd1 vssd1 vccd1 vccd1 _04363_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16981_ _09891_ _10002_ vssd1 vssd1 vccd1 vccd1 _10003_ sky130_fd_sc_hd__nand2_1
XFILLER_27_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18720_ _02822_ rbzero.wall_tracer.rayAddendY\[8\] _02887_ _02917_ vssd1 vssd1 vccd1
+ vccd1 _02918_ sky130_fd_sc_hd__a211o_1
X_15932_ _08516_ _08408_ vssd1 vssd1 vccd1 vccd1 _09027_ sky130_fd_sc_hd__nor2_1
X_11055_ rbzero.tex_b1\[10\] rbzero.tex_b1\[11\] _04325_ vssd1 vssd1 vccd1 vccd1 _04327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15863_ _08696_ _08950_ _08946_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__o21ba_1
X_18651_ _02844_ _02847_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__a21o_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _01891_ _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__xor2_2
X_14814_ rbzero.wall_tracer.stepDistY\[-2\] _07975_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07976_ sky130_fd_sc_hd__mux2_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _08369_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__buf_4
X_18582_ _02786_ _02787_ _02788_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a21o_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_101 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_101/HI zeros[8] sky130_fd_sc_hd__conb_1
XFILLER_205_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_112 vssd1 vssd1 vccd1 vccd1 ones[3] top_ew_algofoogle_112/LO sky130_fd_sc_hd__conb_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_123 vssd1 vssd1 vccd1 vccd1 ones[14] top_ew_algofoogle_123/LO sky130_fd_sc_hd__conb_1
X_17533_ _01823_ _01824_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__nor2_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _07894_ _07909_ _07912_ _07903_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__a211o_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ rbzero.debug_overlay.facingX\[-8\] _05117_ _05122_ rbzero.debug_overlay.facingX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a22o_1
XFILLER_189_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _04248_ vssd1 vssd1 vccd1 vccd1 _04250_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17464_ _08123_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__buf_8
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14676_ _07842_ _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__xnor2_2
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11888_ _04641_ _05053_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or3b_1
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16415_ _09497_ _09505_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__xnor2_1
X_19203_ _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__buf_2
X_13627_ _06682_ _06692_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__xnor2_2
X_17395_ _01672_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__xnor2_1
X_10839_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04203_ vssd1 vssd1 vccd1 vccd1 _04213_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ _09420_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__nand3_1
XFILLER_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19134_ rbzero.spi_registers.new_texadd\[0\]\[19\] _03155_ _03167_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__o211a_1
XFILLER_201_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13558_ _06671_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_160_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19065_ rbzero.spi_registers.new_mapd\[15\] _03120_ _03128_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00772_ sky130_fd_sc_hd__o211a_1
X_12509_ net9 _05642_ _05678_ _05683_ _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a41o_2
X_16277_ _09005_ _08553_ _09273_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__or3_1
XFILLER_121_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13489_ _06512_ _06590_ _06586_ _06554_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__a211o_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _02227_ _02231_ _02233_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a21oi_1
X_15228_ _06034_ _06074_ _08322_ _08158_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__a31o_1
XFILLER_172_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15159_ rbzero.debug_overlay.playerX\[-4\] rbzero.debug_overlay.playerX\[-5\] _08215_
+ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__or3_1
XFILLER_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19967_ rbzero.pov.ready_buffer\[46\] _03438_ _03610_ _03618_ vssd1 vssd1 vccd1 vccd1
+ _03619_ sky130_fd_sc_hd__a211o_1
XFILLER_141_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18918_ rbzero.pov.spi_buffer\[66\] rbzero.pov.ready_buffer\[66\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_68_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19898_ rbzero.debug_overlay.playerX\[-8\] _03565_ vssd1 vssd1 vccd1 vccd1 _03566_
+ sky130_fd_sc_hd__or2_1
XFILLER_110_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18849_ rbzero.pov.spi_buffer\[33\] rbzero.pov.ready_buffer\[33\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21860_ net386 _01449_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20811_ clknet_leaf_58_i_clk _00400_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21791_ net317 _01380_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20742_ rbzero.traced_texVinit\[7\] _09759_ _03937_ _09721_ vssd1 vssd1 vccd1 vccd1
+ _01641_ sky130_fd_sc_hd__a22o_1
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20673_ _03888_ _03890_ _03889_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a21boi_1
XFILLER_51_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20488__335 clknet_1_1__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__inv_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21225_ clknet_leaf_24_i_clk _00814_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21156_ clknet_leaf_12_i_clk _00745_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20107_ rbzero.pov.ready_buffer\[5\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__and3_1
X_21087_ clknet_leaf_97_i_clk _00676_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20038_ rbzero.debug_overlay.facingX\[-2\] _03658_ vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__or2_1
XFILLER_74_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12860_ _06033_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nand2_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ rbzero.tex_r0\[51\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__and3_1
XFILLER_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _05948_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__nand2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ net135 _01578_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _07690_ _07691_ _07699_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__nand3_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__buf_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14461_ _07630_ _07631_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__nand2_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ gpout0.hpos\[8\] _04843_ _04845_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16200_ _08516_ _08429_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__nor2_1
X_13412_ _06512_ _06582_ _06504_ _06498_ _06554_ _06578_ vssd1 vssd1 vccd1 vccd1 _06583_
+ sky130_fd_sc_hd__mux4_1
X_10624_ _04100_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__clkbuf_1
X_17180_ _10182_ _10199_ vssd1 vssd1 vccd1 vccd1 _10200_ sky130_fd_sc_hd__xnor2_1
X_14392_ _07560_ _07562_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _09222_ _09224_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__xnor2_4
XFILLER_10_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13343_ _06482_ _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__or2_1
X_10555_ rbzero.tex_r0\[56\] rbzero.tex_r0\[55\] _04055_ vssd1 vssd1 vccd1 vccd1 _04064_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16062_ _08557_ _09011_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__nand2_1
XFILLER_170_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13274_ _06439_ _06440_ _06442_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__o211a_1
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ rbzero.tex_r1\[22\] rbzero.tex_r1\[23\] _04024_ vssd1 vssd1 vccd1 vccd1 _04026_
+ sky130_fd_sc_hd__mux2_1
X_15013_ _08116_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__clkbuf_4
X_12225_ rbzero.tex_g1\[29\] _04981_ _04831_ _04939_ vssd1 vssd1 vccd1 vccd1 _05412_
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ rbzero.pov.spi_buffer\[48\] rbzero.pov.spi_buffer\[49\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03522_ sky130_fd_sc_hd__mux2_1
X_12156_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _04933_ vssd1 vssd1 vccd1 vccd1 _05344_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ rbzero.tex_b0\[50\] rbzero.tex_b0\[49\] _04351_ vssd1 vssd1 vccd1 vccd1 _04354_
+ sky130_fd_sc_hd__mux2_1
X_19752_ rbzero.pov.spi_buffer\[15\] rbzero.pov.spi_buffer\[16\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux2_1
X_16964_ _09697_ _09699_ vssd1 vssd1 vccd1 vccd1 _09986_ sky130_fd_sc_hd__or2b_1
X_12087_ _05272_ _05274_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__or3_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18703_ _09753_ _02893_ _02894_ _02902_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__a31o_1
X_15915_ _09007_ _09009_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__xnor2_1
X_11038_ rbzero.tex_b1\[18\] rbzero.tex_b1\[19\] _04314_ vssd1 vssd1 vccd1 vccd1 _04318_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16895_ _09915_ _09916_ vssd1 vssd1 vccd1 vccd1 _09917_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _02835_ _02836_ _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a211o_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _08868_ _08900_ _08907_ _08940_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__and4_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _08135_ _02773_ _02774_ _09745_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a31o_1
X_15777_ _08849_ _08848_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__nand2_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12989_ rbzero.wall_tracer.trackDistX\[8\] vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__inv_2
XFILLER_166_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17516_ _01806_ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__nand2_1
X_14728_ _07894_ _07895_ _07896_ _06619_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__o211a_1
XFILLER_178_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18496_ _06082_ _06083_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__nand2_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17447_ _10328_ _10351_ _01739_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14659_ _07333_ _07401_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__and2_1
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17378_ _09146_ _09687_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__and2_1
XFILLER_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19117_ rbzero.spi_registers.texadd0\[11\] _03156_ vssd1 vssd1 vccd1 vccd1 _03159_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16329_ rbzero.wall_tracer.stepDistX\[6\] _09045_ vssd1 vssd1 vccd1 vccd1 _09421_
+ sky130_fd_sc_hd__nand2_2
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19048_ _03084_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__clkbuf_8
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21010_ clknet_leaf_78_i_clk _00599_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19661__42 clknet_1_0__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21912_ net438 _01501_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
X_21843_ net369 _01432_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21774_ net300 _01363_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20725_ _03728_ clknet_1_0__leaf__05820_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and2_2
XFILLER_196_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20656_ _03876_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__a21o_1
XFILLER_108_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20587_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03821_
+ sky130_fd_sc_hd__nor2_1
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__buf_4
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21208_ clknet_leaf_10_i_clk _00797_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21139_ clknet_leaf_23_i_clk _00728_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13961_ _06732_ _06769_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__nor2_1
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700_ _08786_ _08793_ _08794_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__a21o_1
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12912_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__buf_2
X_16680_ _09744_ vssd1 vssd1 vccd1 vccd1 _09751_ sky130_fd_sc_hd__clkbuf_8
X_20542__384 clknet_1_0__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__inv_2
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _07061_ _06885_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__o21ba_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15631_ _08716_ _08723_ _08725_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__a21oi_2
X_12843_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__nor2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20241__112 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__inv_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15562_ _08654_ _08656_ _08629_ _08653_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__o2bb2a_1
X_18350_ _02569_ rbzero.wall_tracer.rayAddendX\[0\] _02568_ vssd1 vssd1 vccd1 vccd1
+ _02584_ sky130_fd_sc_hd__o21a_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12774_ net71 _05944_ _05941_ _05055_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a221o_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _10190_ _10318_ _10319_ vssd1 vssd1 vccd1 vccd1 _10320_ sky130_fd_sc_hd__a21oi_1
X_14513_ _07676_ _07679_ _07681_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__and3_1
XFILLER_15_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _04914_ vssd1 vssd1 vccd1 vccd1 _04915_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _08370_ _08228_ _08586_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__o21ai_1
X_18281_ _05120_ rbzero.wall_tracer.rayAddendX\[-6\] _02520_ vssd1 vssd1 vccd1 vccd1
+ _02521_ sky130_fd_sc_hd__o21ai_1
XFILLER_203_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17232_ _10124_ _10250_ _10251_ vssd1 vssd1 vccd1 vccd1 _10252_ sky130_fd_sc_hd__a21o_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14444_ _07606_ _07613_ _07614_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ rbzero.row_render.size\[6\] _04839_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nor2_1
XFILLER_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ _04091_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17163_ _08338_ _08499_ vssd1 vssd1 vccd1 vccd1 _10183_ sky130_fd_sc_hd__nor2_1
XFILLER_35_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _07491_ _07543_ _07545_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__a21o_1
X_11587_ rbzero.texV\[3\] _04775_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__a21boi_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _09060_ _09062_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__and2b_1
XFILLER_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _06373_ _06377_ _06415_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o21a_1
X_17094_ _10113_ _10114_ vssd1 vssd1 vccd1 vccd1 _10115_ sky130_fd_sc_hd__nor2_1
X_10538_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16045_ _09136_ _09138_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__xnor2_1
X_13257_ _06328_ _06427_ _04444_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10469_ rbzero.tex_r1\[30\] rbzero.tex_r1\[31\] _04013_ vssd1 vssd1 vccd1 vccd1 _04017_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12208_ rbzero.tex_g1\[4\] _04935_ _05305_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13188_ _04443_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nand2_1
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ _03513_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
X_12139_ _04920_ _05322_ _05326_ _04955_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a211o_1
XFILLER_42_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17996_ _08499_ _09621_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__nor2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19735_ rbzero.pov.spi_buffer\[7\] rbzero.pov.spi_buffer\[8\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _06433_ _09691_ _09692_ _09686_ vssd1 vssd1 vccd1 vccd1 _09969_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19666_ clknet_1_1__leaf__03457_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__buf_1
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16878_ _08952_ _09362_ vssd1 vssd1 vccd1 vccd1 _09900_ sky130_fd_sc_hd__nor2_1
XFILLER_93_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18617_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15829_ _08274_ _08473_ _08458_ _08296_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__o22a_1
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19597_ _03427_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18548_ _05132_ rbzero.wall_tracer.rayAddendY\[-4\] vssd1 vssd1 vccd1 vccd1 _02759_
+ sky130_fd_sc_hd__and2_1
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18479_ rbzero.debug_overlay.playerY\[0\] _06130_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02703_ sky130_fd_sc_hd__mux2_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21490_ net208 _01079_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22042_ clknet_leaf_37_i_clk _01631_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21826_ net352 _01415_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21757_ net283 _01346_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _04579_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__or2_1
XFILLER_141_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20708_ _04436_ _08141_ _04437_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__o21ai_1
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12490_ _05661_ _05640_ _05667_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a31o_1
XFILLER_180_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21688_ clknet_leaf_6_i_clk _01277_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _04631_ _04632_ _04422_ _04426_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__o211a_1
XFILLER_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20639_ _03861_ _03862_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nor2_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14160_ _07303_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__buf_2
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ _04549_ _04552_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or2_1
X_13111_ _06078_ _06281_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or2_1
X_14091_ _06718_ _07078_ _06727_ _06540_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__o22a_1
XFILLER_180_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13042_ _06144_ _06113_ rbzero.map_rom.f2 rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1
+ vccd1 _06218_ sky130_fd_sc_hd__or4_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17850_ _09670_ _02007_ _01898_ _09662_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__o22ai_1
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16801_ _06105_ _09828_ _09829_ _09812_ _09830_ vssd1 vssd1 vccd1 vccd1 _09831_ sky130_fd_sc_hd__o311a_1
XFILLER_152_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17781_ _01958_ _01960_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nor2_1
X_14993_ _08106_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19520_ rbzero.spi_registers.new_texadd\[0\]\[2\] _02483_ _03381_ vssd1 vssd1 vccd1
+ vccd1 _03388_ sky130_fd_sc_hd__mux2_1
X_16732_ rbzero.map_rom.f2 _08218_ vssd1 vssd1 vccd1 vccd1 _09770_ sky130_fd_sc_hd__nor2_1
X_13944_ _06742_ _06743_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__nand2_1
XFILLER_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ _04408_ _02930_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__nor3b_4
X_13875_ _06959_ _06857_ _07045_ _06772_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__o22a_1
X_16663_ _04420_ _09739_ _09742_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o21a_1
XFILLER_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18402_ _02626_ _02627_ _02632_ _04434_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__o22a_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15614_ _08363_ _08701_ _08702_ _08704_ _08700_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__a32oi_4
X_12826_ _05999_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__or3_1
XFILLER_62_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19382_ _02483_ rbzero.spi_registers.new_sky\[2\] _03309_ vssd1 vssd1 vccd1 vccd1
+ _03312_ sky130_fd_sc_hd__mux2_1
X_16594_ _09678_ _09683_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__xor2_1
XFILLER_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20553__14 clknet_1_0__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XFILLER_203_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18333_ _02558_ _02561_ _02559_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a21bo_1
X_15545_ _08636_ _08639_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__and2_1
X_12757_ _05932_ _05934_ _05918_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__o21a_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ rbzero.floor_leak\[5\] _04810_ _04887_ rbzero.floor_leak\[4\] _04897_ vssd1
+ vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__o221a_1
X_15476_ _08546_ _08570_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18264_ rbzero.spi_registers.new_texadd\[2\]\[21\] rbzero.spi_registers.spi_buffer\[21\]
+ _02478_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_187_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12688_ _03975_ _04420_ _05822_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__mux2_1
XFILLER_124_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17215_ _10056_ _10111_ _10109_ vssd1 vssd1 vccd1 vccd1 _10235_ sky130_fd_sc_hd__a21oi_1
X_14427_ _07588_ _07595_ _07597_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__a21oi_2
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _04785_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__and2_2
X_18195_ _02176_ _02461_ _02364_ rbzero.wall_tracer.trackDistY\[8\] vssd1 vssd1 vccd1
+ vccd1 _00569_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_156_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17146_ _10060_ _10061_ vssd1 vssd1 vccd1 vccd1 _10166_ sky130_fd_sc_hd__nand2_1
X_14358_ _07527_ _07528_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__nor2_1
XFILLER_156_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03784_ clknet_0__03784_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03784_
+ sky130_fd_sc_hd__clkbuf_16
X_13309_ _06478_ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__xnor2_4
X_17077_ _09969_ _09979_ vssd1 vssd1 vccd1 vccd1 _10098_ sky130_fd_sc_hd__nor2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14289_ _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__nand2_1
XFILLER_171_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16028_ _09117_ _09121_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__nor2_1
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20248__118 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__inv_2
XFILLER_85_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17979_ _02177_ _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__and2_1
X_20226__98 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__inv_2
X_19718_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20990_ clknet_leaf_25_i_clk _00579_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21611_ clknet_leaf_88_i_clk _01200_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21542_ clknet_leaf_71_i_clk _01131_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21473_ net191 _01062_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22025_ clknet_leaf_39_i_clk _01614_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11990_ rbzero.row_render.texu\[4\] _04958_ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_
+ sky130_fd_sc_hd__a21oi_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10941_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _04259_ vssd1 vssd1 vccd1 vccd1 _04267_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ _06717_ _06785_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__or2_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10872_ rbzero.tex_g0\[34\] rbzero.tex_g0\[33\] _04226_ vssd1 vssd1 vccd1 vccd1 _04231_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _05780_ _05763_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nor2_1
X_21809_ net335 _01398_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _06756_ _06761_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__nand2_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _07992_ _08393_ _07996_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__a21o_1
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ net43 _05719_ _05720_ net46 _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a221o_1
XFILLER_129_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ _08328_ _08343_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__nor2_1
XFILLER_40_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20353__213 clknet_1_1__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__inv_2
XFILLER_71_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12473_ _05654_ _05640_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__or2b_1
XFILLER_138_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19689__67 clknet_1_1__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_32_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ _09926_ _10019_ _10020_ vssd1 vssd1 vccd1 vccd1 _10021_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14212_ _07304_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__and2_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11424_ rbzero.spi_registers.texadd0\[1\] _04535_ _04614_ _04615_ _04454_ vssd1 vssd1
+ vccd1 vccd1 _04616_ sky130_fd_sc_hd__o221a_1
X_15192_ _06263_ _08280_ _08286_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__o21ai_4
XANTENNA_8 _07935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14143_ _07304_ _07312_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__xor2_1
XFILLER_193_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11355_ rbzero.spi_registers.texadd1\[20\] _04545_ _04536_ _04546_ vssd1 vssd1 vccd1
+ vccd1 _04547_ sky130_fd_sc_hd__a211o_1
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ _07215_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__xor2_4
X_18951_ _03059_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ rbzero.spi_registers.texadd1\[10\] _04460_ vssd1 vssd1 vccd1 vccd1 _04478_
+ sky130_fd_sc_hd__and2_1
XFILLER_152_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17902_ _10288_ _09433_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nor2_1
XFILLER_117_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13025_ _06197_ rbzero.wall_tracer.trackDistX\[-4\] _06198_ _06200_ vssd1 vssd1 vccd1
+ vccd1 _06201_ sky130_fd_sc_hd__o211ai_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18882_ _02966_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__buf_4
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17833_ _02058_ _02043_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__or2b_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17764_ _02052_ _02053_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14976_ _08097_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19503_ _03378_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__clkbuf_1
X_16715_ rbzero.traced_texa\[7\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a22o_1
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ _06879_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__xnor2_1
X_17695_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__nand2_1
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19434_ _02485_ rbzero.spi_registers.new_other\[3\] _03338_ vssd1 vssd1 vccd1 vccd1
+ _03342_ sky130_fd_sc_hd__mux2_1
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16646_ _09733_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__clkbuf_1
X_13858_ _07025_ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__xor2_1
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ net126 _05946_ _05958_ _05940_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a211oi_2
XFILLER_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19365_ _03212_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__buf_4
X_16577_ _09315_ _09306_ _08369_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__a21oi_2
XFILLER_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13789_ _06959_ _06719_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__or2_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18316_ _02551_ _02552_ _08136_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a21oi_1
X_15528_ _08619_ _08621_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__and2_1
XFILLER_163_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19296_ rbzero.spi_registers.new_texadd\[3\]\[15\] _03254_ _03261_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__o211a_1
XFILLER_37_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18247_ _02498_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15459_ _08304_ _08553_ _08551_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18178_ _02446_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__clkbuf_1
X_17129_ _10058_ _10074_ _10148_ vssd1 vssd1 vccd1 vccd1 _10149_ sky130_fd_sc_hd__a21bo_1
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20140_ _03728_ _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__and3_1
Xclkbuf_0__03798_ _03798_ vssd1 vssd1 vccd1 vccd1 clknet_0__03798_ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ rbzero.pov.ready_buffer\[32\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__and3_1
XFILLER_135_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_1_i_clk clknet_1_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0_1_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20973_ clknet_leaf_61_i_clk _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20302__167 clknet_1_0__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__inv_2
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21525_ clknet_leaf_84_i_clk _01114_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21456_ net174 _01045_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21387_ clknet_leaf_8_i_clk _00976_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ rbzero.tex_b0\[34\] rbzero.tex_b0\[33\] _04362_ vssd1 vssd1 vccd1 vccd1 _04371_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 o_gpout[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__buf_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11071_ rbzero.tex_b1\[2\] rbzero.tex_b1\[3\] _04325_ vssd1 vssd1 vccd1 vccd1 _04335_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22008_ net130 _01597_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _07989_ _07921_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__and2_1
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11973_ _05157_ _05159_ _05161_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__or3_1
X_14761_ _07894_ _07926_ _07927_ _07903_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__a211o_1
XFILLER_99_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16500_ _09463_ _09589_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__03787_ clknet_0__03787_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03787_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10924_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _04248_ vssd1 vssd1 vccd1 vccd1 _04258_
+ sky130_fd_sc_hd__mux2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06826_ _06827_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__and2b_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17480_ _01672_ _01687_ _01685_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a21o_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _07067_ _07826_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__nand2_1
XFILLER_189_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _08166_ _08666_ vssd1 vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__or2_1
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ rbzero.tex_g0\[42\] rbzero.tex_g0\[41\] _04215_ vssd1 vssd1 vccd1 vccd1 _04222_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _06804_ _06811_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__nand2_1
XFILLER_198_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19150_ rbzero.spi_registers.texadd1\[1\] _03176_ vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__or2_1
X_16362_ _09452_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__nor2_1
X_13574_ _06707_ _06741_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__nand2_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _04185_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__clkbuf_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__or2_1
XFILLER_158_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15313_ _08161_ _08404_ _08406_ _08407_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__o211a_2
X_12525_ _05704_ _05297_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nand2_1
X_16293_ _09280_ _09282_ _09284_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__o21ai_1
X_19081_ rbzero.mapdxw\[1\] _03121_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__or2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18032_ _02248_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20568__4 clknet_1_1__leaf__03457_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
X_15244_ _06076_ _08158_ _08320_ _08338_ _08069_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__o32a_1
X_12456_ net7 net6 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__nor2_2
XFILLER_138_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ _04575_ _04594_ _04596_ _04598_ _04452_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__o221a_1
X_15175_ _07933_ _07934_ _08143_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__a21o_1
X_12387_ rbzero.tex_b1\[34\] _04914_ _04981_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a21o_1
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14126_ _07280_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__nor2_1
XFILLER_119_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _04525_ _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__nor2_1
XFILLER_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19983_ _03212_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__buf_4
XFILLER_180_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18934_ rbzero.spi_registers.spi_counter\[4\] rbzero.spi_registers.spi_counter\[3\]
+ rbzero.spi_registers.spi_counter\[2\] _02945_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor4_1
X_14057_ _06640_ _06719_ _07225_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__o21a_1
X_11269_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__clkbuf_4
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13008_ rbzero.wall_tracer.trackDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__inv_2
X_18865_ _03013_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
X_17816_ _08814_ _10093_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__nor2_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18796_ rbzero.pov.spi_buffer\[8\] rbzero.pov.ready_buffer\[8\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02977_ sky130_fd_sc_hd__mux2_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17747_ _01842_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14959_ _08065_ _08086_ _08087_ _08085_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__o211a_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17678_ _01769_ _01967_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__or2_1
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19417_ _03332_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16629_ _09717_ _09718_ vssd1 vssd1 vccd1 vccd1 _09719_ sky130_fd_sc_hd__or2_2
XFILLER_189_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19348_ rbzero.spi_registers.new_floor\[1\] rbzero.spi_registers.got_new_floor _03097_
+ _04409_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a31o_1
XFILLER_176_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19279_ _03212_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_149_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21310_ clknet_leaf_35_i_clk _00899_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19668__48 clknet_1_0__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21241_ clknet_leaf_6_i_clk _00830_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21172_ clknet_leaf_14_i_clk _00761_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20123_ _05648_ _05651_ _03091_ _04657_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and4b_1
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20054_ rbzero.debug_overlay.facingY\[-6\] _03676_ _03678_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01211_ sky130_fd_sc_hd__a211o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20956_ clknet_leaf_63_i_clk _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ clknet_leaf_46_i_clk _00476_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _04108_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _04072_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12310_ _04946_ _05493_ _05494_ _05495_ _04952_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__o221a_1
XFILLER_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21508_ clknet_leaf_82_i_clk _01097_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _06405_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__xnor2_2
XFILLER_155_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ rbzero.tex_g1\[62\] _04830_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__or2_1
X_21439_ net157 _01028_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12172_ _04920_ _05355_ _05359_ _04903_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a211o_1
X_11123_ _04214_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__clkbuf_4
X_20465__314 clknet_1_0__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__inv_2
X_16980_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10002_ sky130_fd_sc_hd__xor2_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _04326_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
X_15931_ _08432_ _08435_ _08430_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__a21bo_1
XFILLER_150_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18650_ _02794_ _05132_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _08616_ _08461_ _08945_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__or3b_1
XFILLER_190_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17601_ _09520_ _09890_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__and2_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14813_ _06670_ _07973_ _07974_ _06516_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__a211o_4
XFILLER_114_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18581_ _02786_ _02787_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__nand3_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _08880_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__o21ai_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_102 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_102/HI zeros[9] sky130_fd_sc_hd__conb_1
XFILLER_188_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17532_ _01820_ _01822_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_79_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_113 vssd1 vssd1 vccd1 vccd1 ones[4] top_ew_algofoogle_113/LO sky130_fd_sc_hd__conb_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _06577_ _07911_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__and2_1
Xtop_ew_algofoogle_124 vssd1 vssd1 vccd1 vccd1 ones[15] top_ew_algofoogle_124/LO sky130_fd_sc_hd__conb_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _04657_ _04651_ _05126_ _05136_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a41o_1
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17463_ _10248_ _10253_ _10369_ _10371_ _01755_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a41o_1
X_10907_ _04249_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14675_ _07830_ _07843_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__a21oi_2
X_11887_ _05066_ _05070_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__or2_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19202_ rbzero.spi_registers.got_new_texadd\[2\] _03100_ vssd1 vssd1 vccd1 vccd1
+ _03207_ sky130_fd_sc_hd__and2_2
X_16414_ _09503_ _09504_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__nor2_1
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10838_ _04212_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__clkbuf_1
X_13626_ _06788_ _06796_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__xnor2_1
X_17394_ _01685_ _01686_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__nor2_1
XFILLER_38_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19133_ rbzero.spi_registers.texadd0\[19\] _03156_ vssd1 vssd1 vccd1 vccd1 _03167_
+ sky130_fd_sc_hd__or2_1
X_16345_ _09430_ _09431_ _09435_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__a21o_1
X_10769_ _04176_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__clkbuf_1
X_13557_ _06686_ _06684_ _06683_ _06469_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19064_ rbzero.map_overlay.i_mapdx\[5\] _03122_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__or2_1
X_12508_ _05686_ _05687_ _05689_ _05665_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__o31a_2
X_16276_ _09248_ _09249_ _09251_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__a21bo_1
XFILLER_160_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13488_ _06508_ _06578_ _06587_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__a21o_1
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18015_ _02225_ _02239_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__or2b_1
XFILLER_201_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12439_ _04940_ _05619_ _05623_ _04812_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a211o_1
XFILLER_161_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15227_ _08320_ _08321_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_17_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ _08252_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__buf_2
XFILLER_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _07236_ _07258_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__o21ai_1
XFILLER_102_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20331__193 clknet_1_0__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__inv_2
X_19966_ _08204_ _03570_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nor2_1
X_15089_ _06341_ _08183_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__nor2_1
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18917_ _03040_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19897_ net40 _03557_ _03095_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__o21a_2
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18848_ _03004_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18779_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__buf_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20810_ clknet_leaf_51_i_clk _00399_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_21790_ net316 _01379_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20741_ rbzero.traced_texVinit\[6\] _09759_ _03937_ _09593_ vssd1 vssd1 vccd1 vccd1
+ _01640_ sky130_fd_sc_hd__a22o_1
XFILLER_169_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20672_ _09732_ _03891_ _03892_ _03740_ rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1
+ _01615_ sky130_fd_sc_hd__a32o_1
XFILLER_17_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20414__268 clknet_1_1__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__inv_2
XFILLER_152_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21224_ clknet_leaf_24_i_clk _00813_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21155_ clknet_leaf_6_i_clk _00744_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20106_ rbzero.debug_overlay.vplaneY\[-5\] _03655_ _03707_ _03695_ vssd1 vssd1 vccd1
+ vccd1 _01234_ sky130_fd_sc_hd__a211o_1
XFILLER_63_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21086_ clknet_leaf_85_i_clk _00675_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20037_ rbzero.debug_overlay.facingX\[-3\] _03663_ _03668_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01203_ sky130_fd_sc_hd__a211o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20308__173 clknet_1_1__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__inv_2
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _04914_ vssd1 vssd1 vccd1 vccd1 _05000_
+ sky130_fd_sc_hd__mux2_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05652_ _05653_ net34 vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__mux2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21988_ net134 _01577_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _04893_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__buf_4
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ clknet_leaf_56_i_clk _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14460_ _07581_ _07629_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__or2_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _04418_ _04847_ _04844_ gpout0.hpos\[7\] _04861_ vssd1 vssd1 vccd1 vccd1
+ _04862_ sky130_fd_sc_hd__o221a_1
XFILLER_183_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ rbzero.tex_r0\[24\] rbzero.tex_r0\[23\] _04099_ vssd1 vssd1 vccd1 vccd1 _04100_
+ sky130_fd_sc_hd__mux2_1
X_13411_ _06501_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__inv_2
XFILLER_186_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14391_ _07507_ _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__nand2_1
XFILLER_70_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _08625_ _09092_ _09223_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__a21oi_4
XFILLER_127_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13342_ _06474_ _06508_ _06510_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__or4_1
X_10554_ _04063_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16061_ _09153_ _09154_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__xnor2_1
X_13273_ _06415_ _06438_ _06441_ _06443_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a211o_1
X_10485_ _04025_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19647__29 clknet_1_1__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_108_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12224_ rbzero.tex_g1\[31\] _05305_ _05410_ _04912_ vssd1 vssd1 vccd1 vccd1 _05411_
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15012_ _03974_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__buf_4
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _03521_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _05339_ _05342_ _04941_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__mux2_1
XFILLER_2_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _04353_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19751_ _03485_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16963_ _09964_ _09984_ vssd1 vssd1 vccd1 vccd1 _09985_ sky130_fd_sc_hd__xnor2_2
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12086_ _04651_ _04419_ _04411_ _04648_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_150_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18702_ _08135_ _02900_ _02901_ _09751_ rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a32o_1
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ _09008_ _08553_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__nor2_1
X_11037_ _04317_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16894_ _09146_ _09131_ vssd1 vssd1 vccd1 vccd1 _09916_ sky130_fd_sc_hd__nor2_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18633_ _02833_ _02834_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__o211ai_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _08909_ _08939_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__nor2_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ rbzero.debug_overlay.vplaneY\[-7\] _02764_ vssd1 vssd1 vccd1 vccd1 _02774_
+ sky130_fd_sc_hd__nand2_1
XFILLER_40_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _08851_ _08853_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__xnor2_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12988_ rbzero.wall_tracer.trackDistX\[10\] vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__inv_2
X_17515_ _01725_ _01717_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__or2b_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14727_ _06540_ _06577_ _07855_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__or3b_1
X_11939_ rbzero.debug_overlay.vplaneY\[-1\] _05108_ _05115_ rbzero.debug_overlay.vplaneY\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a22o_1
X_18495_ _02715_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17446_ _10348_ _10350_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__and2b_1
X_14658_ _06758_ _06738_ _07331_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__a21oi_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _06774_ _06778_ _06777_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__a21oi_1
X_17377_ _01668_ _01669_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__xor2_1
X_14589_ _07045_ _07476_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__nor2_1
XFILLER_158_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19116_ rbzero.spi_registers.new_texadd\[0\]\[10\] _03155_ _03157_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__o211a_1
XFILLER_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16328_ _09416_ _09419_ vssd1 vssd1 vccd1 vccd1 _09420_ sky130_fd_sc_hd__xor2_1
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ rbzero.spi_registers.got_new_vinf _03100_ rbzero.row_render.vinf vssd1 vssd1
+ vccd1 vccd1 _03117_ sky130_fd_sc_hd__a21o_1
X_16259_ _09350_ _09351_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__nor2_1
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19949_ _03556_ _03604_ _03565_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__o21a_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21911_ net437 _01500_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21842_ net368 _01431_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21773_ net299 _01362_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20494__340 clknet_1_1__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__inv_2
X_20724_ _03932_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__buf_1
XFILLER_208_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20655_ _03871_ _03875_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__nand2_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20586_ _03816_ _03817_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__and2_1
XFILLER_192_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20338__199 clknet_1_1__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__inv_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21207_ clknet_leaf_10_i_clk _00796_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21138_ clknet_leaf_21_i_clk _00727_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21069_ clknet_leaf_83_i_clk _00658_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13960_ _07075_ _07083_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__and2_1
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12911_ _06076_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__inv_2
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13891_ _06875_ _06851_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__and2b_1
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15630_ _08700_ _08724_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__or2_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _06002_ _06009_ _06010_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__or4bb_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _08367_ _08655_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__and2_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ net49 _05945_ _05947_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a211o_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17300_ _09528_ _09186_ _09669_ _08814_ vssd1 vssd1 vccd1 vccd1 _10319_ sky130_fd_sc_hd__o22a_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14512_ _07648_ _07662_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__xnor2_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__clkbuf_8
X_18280_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] _02519_
+ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a21o_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _08370_ _08228_ _08586_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__or3_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _10017_ _10003_ _10121_ vssd1 vssd1 vccd1 vccd1 _10251_ sky130_fd_sc_hd__and3_1
XFILLER_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14443_ _07608_ _07612_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__nor2_1
X_11655_ gpout0.hpos\[7\] _04844_ _04843_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1
+ _04845_ sky130_fd_sc_hd__a22o_1
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ rbzero.tex_r0\[32\] rbzero.tex_r0\[31\] _04088_ vssd1 vssd1 vccd1 vccd1 _04091_
+ sky130_fd_sc_hd__mux2_1
X_17162_ _10078_ _10086_ _10181_ vssd1 vssd1 vccd1 vccd1 _10182_ sky130_fd_sc_hd__a21oi_1
XFILLER_161_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _04776_ sky130_fd_sc_hd__nand2_1
XFILLER_35_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14374_ _07306_ _07361_ _07489_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__o21a_1
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ _09175_ _09206_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__xnor2_2
XFILLER_127_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10537_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__buf_4
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13325_ _04444_ _06366_ _06368_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__a21o_1
X_17093_ _09992_ _10024_ _10112_ vssd1 vssd1 vccd1 vccd1 _10114_ sky130_fd_sc_hd__and3_1
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _09078_ _09137_ vssd1 vssd1 vccd1 vccd1 _09138_ sky130_fd_sc_hd__nor2_1
X_10468_ _04016_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__clkbuf_1
X_13256_ rbzero.wall_tracer.visualWallDist\[9\] _04428_ vssd1 vssd1 vccd1 vccd1 _06427_
+ sky130_fd_sc_hd__or2_1
X_12207_ rbzero.tex_g1\[5\] _04981_ _04831_ _04939_ vssd1 vssd1 vccd1 vccd1 _05394_
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13187_ _06308_ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__xnor2_1
X_10399_ _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__clkbuf_4
XFILLER_151_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ _05191_ _05323_ _05324_ _05325_ _04937_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__o221a_1
X_19803_ rbzero.pov.spi_buffer\[39\] rbzero.pov.spi_buffer\[40\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03513_ sky130_fd_sc_hd__mux2_1
X_17995_ _02124_ _02216_ _02219_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__o21a_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16946_ _09965_ _09967_ vssd1 vssd1 vccd1 vccd1 _09968_ sky130_fd_sc_hd__xor2_2
X_12069_ rbzero.tex_r1\[51\] _04924_ _05257_ _04944_ vssd1 vssd1 vccd1 vccd1 _05258_
+ sky130_fd_sc_hd__o211a_1
X_19734_ _03476_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16877_ _09660_ _09643_ vssd1 vssd1 vccd1 vccd1 _09899_ sky130_fd_sc_hd__or2b_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18616_ _05127_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__buf_2
XFILLER_93_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20443__294 clknet_1_1__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__inv_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _08922_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__inv_2
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19596_ rbzero.spi_registers.new_texadd\[1\]\[15\] rbzero.spi_registers.spi_buffer\[15\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18547_ _05132_ rbzero.wall_tracer.rayAddendY\[-4\] vssd1 vssd1 vccd1 vccd1 _02758_
+ sky130_fd_sc_hd__nor2_1
X_15759_ _08843_ _08845_ _08850_ _08851_ _08853_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__a32o_1
X_18478_ _02702_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17429_ _01720_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__xor2_1
XFILLER_53_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22041_ clknet_leaf_34_i_clk _01630_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20526__369 clknet_1_1__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__inv_2
XFILLER_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21825_ net351 _01414_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21756_ net282 _01345_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20707_ rbzero.texV\[10\] _03814_ _03819_ _03921_ vssd1 vssd1 vccd1 vccd1 _01621_
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21687_ clknet_leaf_6_i_clk _01276_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _04628_ _04589_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__nor2_1
XFILLER_196_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20638_ rbzero.texV\[-1\] _03814_ _03819_ _03863_ vssd1 vssd1 vccd1 vccd1 _01610_
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ _03970_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nand2_1
X_20271__139 clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__inv_2
XFILLER_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13110_ _06078_ _06281_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
XFILLER_192_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ _07260_ _07221_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__nand2_1
XFILLER_30_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13041_ _06163_ _06215_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__a21o_4
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20546__7 clknet_1_1__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16800_ _09822_ _09111_ vssd1 vssd1 vccd1 vccd1 _09830_ sky130_fd_sc_hd__nand2_1
X_17780_ _01994_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14992_ rbzero.wall_tracer.stepDistX\[1\] _07996_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08106_ sky130_fd_sc_hd__mux2_1
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16731_ rbzero.map_rom.f2 _08218_ vssd1 vssd1 vccd1 vccd1 _09769_ sky130_fd_sc_hd__and2_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13943_ _07073_ _07084_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a21bo_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19450_ rbzero.spi_registers.spi_done _02475_ _02476_ vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__and3_1
X_16662_ _04420_ _09739_ _09730_ vssd1 vssd1 vccd1 vccd1 _09742_ sky130_fd_sc_hd__a21oi_1
X_13874_ _06798_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__clkbuf_4
X_18401_ _02614_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__xnor2_1
X_15613_ _08661_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__xnor2_2
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12825_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__nor2_1
X_19381_ _03311_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
X_16593_ _09679_ _09681_ _09682_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__o21a_1
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18332_ _02557_ _02562_ _02563_ _02567_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a31o_1
X_15544_ _08178_ _08439_ _08636_ _08638_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__or4bb_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12756_ net44 _05910_ _05909_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__a31o_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11707_ rbzero.floor_leak\[3\] _04889_ _04886_ rbzero.floor_leak\[4\] _04896_ vssd1
+ vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18263_ _02506_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15475_ _08568_ _08569_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__nand2_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12687_ _03969_ _04575_ _04452_ _04628_ _05822_ net23 vssd1 vssd1 vccd1 vccd1 _05866_
+ sky130_fd_sc_hd__mux4_1
XFILLER_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17214_ _10179_ _10233_ vssd1 vssd1 vccd1 vccd1 _10234_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14426_ _07478_ _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__or2_1
X_11638_ _04781_ _04784_ _04806_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a21oi_4
X_18194_ _02459_ _02460_ _02337_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__o21a_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17145_ _10163_ _10164_ vssd1 vssd1 vccd1 vccd1 _10165_ sky130_fd_sc_hd__xor2_1
XFILLER_156_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19703__80 clknet_1_0__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
X_14357_ _07472_ _07526_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03783_ clknet_0__03783_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03783_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11569_ rbzero.texV\[6\] _04757_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nand3_1
X_13308_ _06356_ _06392_ _06415_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__o21a_2
X_17076_ _10091_ _10096_ vssd1 vssd1 vccd1 vccd1 _10097_ sky130_fd_sc_hd__xnor2_1
X_14288_ _07415_ _07441_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__xor2_1
XFILLER_170_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16027_ _09117_ _09121_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__and2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13239_ rbzero.wall_tracer.visualWallDist\[10\] _04428_ vssd1 vssd1 vccd1 vccd1 _06410_
+ sky130_fd_sc_hd__or2_1
XFILLER_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17978_ _02178_ _02180_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__nand2_1
XFILLER_85_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16929_ _09949_ _09950_ vssd1 vssd1 vccd1 vccd1 _09951_ sky130_fd_sc_hd__and2b_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19717_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19579_ rbzero.spi_registers.new_texadd\[1\]\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21610_ clknet_leaf_89_i_clk _01199_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21541_ clknet_leaf_71_i_clk _01130_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21472_ net190 _01061_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20423_ clknet_1_0__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__buf_1
XFILLER_88_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22024_ clknet_leaf_55_i_clk _01613_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _04266_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _04230_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ net19 net18 vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__nor2_1
X_21808_ net334 _01397_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _06757_ _06758_ _06756_ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nand4_1
XFILLER_197_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12541_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__inv_2
X_21739_ net265 _01328_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_i_clk clknet_1_1_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _08345_ _08347_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12472_ _05650_ _05651_ _05652_ _05653_ _05646_ net7 vssd1 vssd1 vccd1 vccd1 _05654_
+ sky130_fd_sc_hd__mux4_1
X_14211_ _07067_ _06741_ _07331_ _07344_ _07381_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__a311o_1
XFILLER_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11423_ rbzero.spi_registers.texadd1\[1\] _04545_ _04536_ vssd1 vssd1 vccd1 vccd1
+ _04615_ sky130_fd_sc_hd__a21o_1
X_15191_ _08284_ _08285_ _08158_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__mux2_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 _07971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11354_ rbzero.spi_registers.texadd3\[20\] _04526_ _04537_ rbzero.spi_registers.texadd2\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a22o_1
X_14142_ _07304_ _07312_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__or2b_1
XFILLER_137_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14073_ _07242_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nor2_2
X_11285_ rbzero.texu_hot\[5\] _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__nand2_1
X_18950_ rbzero.spi_registers.spi_buffer\[6\] _02489_ _03052_ vssd1 vssd1 vccd1 vccd1
+ _03059_ sky130_fd_sc_hd__mux2_1
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17901_ _01697_ _10214_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__nor2_1
X_13024_ rbzero.wall_tracer.trackDistX\[1\] _06199_ rbzero.wall_tracer.trackDistX\[-3\]
+ _06180_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__o22a_1
X_18881_ _03021_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17832_ _02005_ _02023_ _02021_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a21o_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _01818_ _09560_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__nor2_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14975_ rbzero.wall_tracer.stepDistX\[-7\] _07935_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08097_ sky130_fd_sc_hd__mux2_1
XFILLER_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16714_ rbzero.traced_texa\[6\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a22o_1
X_19502_ rbzero.spi_registers.new_mapd\[15\] rbzero.spi_registers.spi_buffer\[15\]
+ _03361_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux2_1
XFILLER_48_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13926_ _07088_ _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17694_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__nor2_1
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19433_ _03341_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ _04447_ _04448_ _09732_ vssd1 vssd1 vccd1 vccd1 _09733_ sky130_fd_sc_hd__and3_1
X_13857_ _06982_ _06731_ _07026_ _07027_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__o22ai_2
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12808_ _05952_ _05949_ gpout5.clk_div\[1\] _05984_ vssd1 vssd1 vccd1 vccd1 _05985_
+ sky130_fd_sc_hd__a31o_1
X_19364_ rbzero.spi_registers.vshift\[2\] _03298_ vssd1 vssd1 vccd1 vccd1 _03301_
+ sky130_fd_sc_hd__or2_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16576_ _09545_ _09555_ _09665_ vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__a21bo_1
XFILLER_16_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13788_ _06790_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _02547_ _02548_ _02550_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__o21ai_1
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15527_ _08619_ _08621_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__nor2_1
XFILLER_176_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12739_ _05888_ _05881_ _05884_ _05889_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and4_1
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19295_ rbzero.spi_registers.texadd3\[15\] _03255_ vssd1 vssd1 vccd1 vccd1 _03261_
+ sky130_fd_sc_hd__or2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18246_ rbzero.spi_registers.new_texadd\[2\]\[12\] rbzero.spi_registers.spi_buffer\[12\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
X_15458_ _08541_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14409_ _07551_ _07574_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__xnor2_1
X_18177_ rbzero.wall_tracer.trackDistY\[6\] _02445_ _02339_ vssd1 vssd1 vccd1 vccd1
+ _02446_ sky130_fd_sc_hd__mux2_1
XFILLER_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _08039_ _08161_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__nor2_2
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17128_ _10075_ _10057_ vssd1 vssd1 vccd1 vccd1 _10148_ sky130_fd_sc_hd__or2b_1
XFILLER_117_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17059_ _08910_ _09680_ vssd1 vssd1 vccd1 vccd1 _10080_ sky130_fd_sc_hd__nor2b_1
XFILLER_144_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03797_ _03797_ vssd1 vssd1 vccd1 vccd1 clknet_0__03797_ sky130_fd_sc_hd__clkbuf_16
XFILLER_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20070_ rbzero.debug_overlay.facingY\[0\] _03676_ _03688_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01217_ sky130_fd_sc_hd__a211o_1
XFILLER_83_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20972_ clknet_leaf_58_i_clk _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21524_ clknet_leaf_84_i_clk _01113_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21455_ net173 _01044_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21386_ clknet_leaf_8_i_clk _00975_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__clkbuf_1
X_11070_ _04334_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
X_20268_ clknet_1_1__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__buf_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__buf_2
XFILLER_103_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22007_ net129 _01596_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ _03766_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _07894_ _07900_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__nor2_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11972_ rbzero.debug_overlay.playerX\[-2\] _05107_ _05113_ rbzero.debug_overlay.playerX\[-4\]
+ _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a221o_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03786_ clknet_0__03786_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03786_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13711_ _06879_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__nor2_1
XFILLER_17_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10923_ _04257_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14691_ _07822_ _07856_ _07861_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a21boi_2
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16430_ _08152_ _09519_ _09520_ _08166_ vssd1 vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__o22ai_1
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _06751_ _06746_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__xor2_1
X_10854_ _04221_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _09288_ _09328_ _09326_ vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__a21oi_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _06742_ _06743_ _06732_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__a21oi_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ rbzero.tex_g1\[10\] rbzero.tex_g1\[11\] _04177_ vssd1 vssd1 vccd1 vccd1 _04185_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20277__145 clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__inv_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _02379_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__clkbuf_1
X_15312_ rbzero.wall_tracer.stepDistX\[-1\] _08357_ vssd1 vssd1 vccd1 vccd1 _08407_
+ sky130_fd_sc_hd__nand2_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19080_ rbzero.spi_registers.new_mapd\[2\] _03119_ _03136_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00779_ sky130_fd_sc_hd__o211a_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _05382_ _05470_ _05551_ _05632_ _05704_ net13 vssd1 vssd1 vccd1 vccd1 _05705_
+ sky130_fd_sc_hd__mux4_1
X_16292_ _09359_ _09383_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18031_ _02301_ _02317_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15243_ _08161_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__clkbuf_8
XFILLER_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12455_ net5 net4 vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__nor2_1
XFILLER_166_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ _03970_ _04597_ _04449_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a21o_1
XFILLER_172_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ rbzero.wall_tracer.stepDistX\[-7\] _06262_ vssd1 vssd1 vccd1 vccd1 _08269_
+ sky130_fd_sc_hd__nor2_1
X_12386_ rbzero.tex_b1\[35\] _04926_ _04928_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__and3_1
XFILLER_197_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ _07288_ _07295_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ rbzero.spi_registers.texadd0\[16\] _04467_ _04528_ vssd1 vssd1 vccd1 vccd1
+ _04529_ sky130_fd_sc_hd__o21ai_1
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19982_ rbzero.pov.ready_buffer\[51\] _03570_ _03610_ _03628_ vssd1 vssd1 vccd1 vccd1
+ _03629_ sky130_fd_sc_hd__a211o_1
XFILLER_180_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18933_ _03048_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
X_14056_ _07135_ _07225_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__or3_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _04459_ rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_2
XFILLER_95_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13007_ rbzero.wall_tracer.trackDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__inv_2
X_11199_ rbzero.tex_b0\[6\] rbzero.tex_b0\[5\] _04395_ vssd1 vssd1 vccd1 vccd1 _04402_
+ sky130_fd_sc_hd__mux2_1
X_18864_ rbzero.pov.spi_buffer\[40\] rbzero.pov.ready_buffer\[40\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17815_ _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__and2_1
X_18795_ _02976_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17746_ _02034_ _02035_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__and2_1
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ rbzero.wall_tracer.visualWallDist\[8\] _08046_ vssd1 vssd1 vccd1 vccd1 _08087_
+ sky130_fd_sc_hd__or2_1
XFILLER_208_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _06748_ _06721_ _06758_ _07079_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__a31o_1
X_17677_ _01769_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__nand2_1
XFILLER_39_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14889_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.trackDistX\[-11\]
+ _08037_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__mux2_1
XFILLER_51_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16628_ _09714_ _09716_ vssd1 vssd1 vccd1 vccd1 _09718_ sky130_fd_sc_hd__and2_1
X_19416_ _02483_ rbzero.spi_registers.new_leak\[2\] _03329_ vssd1 vssd1 vccd1 vccd1
+ _03332_ sky130_fd_sc_hd__mux2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16559_ _09646_ _09648_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__nand2_1
X_19347_ rbzero.spi_registers.new_floor\[0\] _03289_ _03291_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00891_ sky130_fd_sc_hd__o211a_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19278_ rbzero.spi_registers.texadd3\[8\] _03242_ vssd1 vssd1 vccd1 vccd1 _03251_
+ sky130_fd_sc_hd__or2_1
XFILLER_206_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18229_ _02488_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21240_ clknet_leaf_24_i_clk _00829_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21171_ clknet_leaf_14_i_clk _00760_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20122_ _04687_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__inv_2
XFILLER_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20053_ rbzero.pov.ready_buffer\[25\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__and3_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ clknet_leaf_65_i_clk _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ clknet_leaf_46_i_clk _00475_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _04066_ vssd1 vssd1 vccd1 vccd1 _04072_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21507_ clknet_leaf_83_i_clk _01096_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ rbzero.tex_g1\[48\] _04905_ _05305_ _05425_ _05426_ vssd1 vssd1 vccd1 vccd1
+ _05427_ sky130_fd_sc_hd__a311o_1
X_21438_ net156 _01027_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _05191_ _05356_ _05357_ _05358_ _04937_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__o221a_1
X_21369_ clknet_leaf_13_i_clk _00958_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11122_ _04361_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15930_ _08377_ _08385_ _08387_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__a21bo_1
X_11053_ rbzero.tex_b1\[11\] rbzero.tex_b1\[12\] _04325_ vssd1 vssd1 vccd1 vccd1 _04326_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _08951_ _08955_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _01889_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__xor2_2
XFILLER_40_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14812_ _06574_ _07881_ _07888_ _06655_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__o211a_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _02776_ _02779_ _02777_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a21bo_1
X_15792_ _08871_ _08886_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__xnor2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _01820_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__nor2_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_103 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_103/HI zeros[10]
+ sky130_fd_sc_hd__conb_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _07806_ _07804_ _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__a21oi_1
Xtop_ew_algofoogle_114 vssd1 vssd1 vccd1 vccd1 ones[5] top_ew_algofoogle_114/LO sky130_fd_sc_hd__conb_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _04731_ _04654_ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__nor3_1
XFILLER_189_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20570__6 clknet_1_1__leaf__03457_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _10246_ _10369_ _10370_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ rbzero.tex_g0\[18\] rbzero.tex_g0\[17\] _04248_ vssd1 vssd1 vccd1 vccd1 _04249_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _07830_ _07843_ _07831_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ _04424_ _04636_ _05074_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a21oi_4
X_16413_ _09388_ _09390_ _09502_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__and3_1
X_19201_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__clkbuf_4
X_13625_ _06789_ _06794_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a21boi_1
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17393_ _01683_ _01684_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__and2_1
X_10837_ rbzero.tex_g0\[50\] rbzero.tex_g0\[49\] _04203_ vssd1 vssd1 vccd1 vccd1 _04212_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19132_ rbzero.spi_registers.new_texadd\[0\]\[18\] _03155_ _03166_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__o211a_1
X_16344_ _09430_ _09431_ _09435_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__nand3_1
XFILLER_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13556_ _06640_ _06708_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__xnor2_4
XFILLER_199_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10768_ rbzero.tex_g1\[18\] rbzero.tex_g1\[19\] _04166_ vssd1 vssd1 vccd1 vccd1 _04176_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19063_ rbzero.spi_registers.new_mapd\[14\] _03120_ _03127_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00771_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_12507_ gpout0.clk_div\[1\] _05638_ _05663_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_
+ sky130_fd_sc_hd__a31o_2
X_16275_ _09244_ _09364_ _09366_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _06633_ _06650_ _06654_ _06655_ _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a32o_4
XFILLER_201_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10699_ _04139_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__clkbuf_1
X_18014_ _02299_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__xnor2_1
X_15226_ rbzero.debug_overlay.playerY\[-2\] _08281_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__o21ai_1
X_12438_ _04827_ _05620_ _05622_ _04918_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__o211a_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15157_ _08250_ _08251_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__or2b_1
XFILLER_126_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12369_ _04818_ _05036_ _05177_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14108_ _07276_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19965_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__clkbuf_4
X_15088_ _06396_ _06397_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__nor2_1
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18916_ rbzero.pov.spi_buffer\[65\] rbzero.pov.ready_buffer\[65\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
X_14039_ _07206_ _07209_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor2_1
XFILLER_80_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03465_ clknet_0__03465_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03465_
+ sky130_fd_sc_hd__clkbuf_16
X_19896_ _08186_ rbzero.pov.ready_buffer\[60\] _03561_ vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18847_ rbzero.pov.spi_buffer\[32\] rbzero.pov.ready_buffer\[32\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18778_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__buf_4
XFILLER_208_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17729_ _02006_ _02018_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20740_ rbzero.traced_texVinit\[5\] _09759_ _03937_ _09868_ vssd1 vssd1 vccd1 vccd1
+ _01639_ sky130_fd_sc_hd__a22o_1
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20671_ _03888_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nand3_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21223_ clknet_leaf_28_i_clk _00812_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21154_ clknet_leaf_6_i_clk _00743_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20105_ rbzero.pov.ready_buffer\[4\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__and3_1
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21085_ clknet_leaf_88_i_clk _00674_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20036_ _04409_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21987_ net133 _01576_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ rbzero.tex_r0\[3\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and3_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ clknet_leaf_48_i_clk _00527_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _04411_ _04849_ _04847_ _04418_ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a221o_1
X_20869_ clknet_leaf_36_i_clk _00458_ vssd1 vssd1 vccd1 vccd1 reg_rgb\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13410_ _06469_ _06568_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__nand2_4
X_10622_ _04054_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14390_ _06757_ _06785_ _07366_ _07309_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__or4b_1
XFILLER_169_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _06385_ _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__xnor2_4
X_10553_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _04055_ vssd1 vssd1 vccd1 vccd1 _04063_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16060_ _08235_ _08340_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__nor2_1
X_13272_ _06414_ _06421_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and2_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ rbzero.tex_r1\[23\] rbzero.tex_r1\[24\] _04024_ vssd1 vssd1 vccd1 vccd1 _04025_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _08115_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12223_ rbzero.tex_g1\[30\] _05236_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__or2_1
XFILLER_68_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20389__246 clknet_1_0__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__inv_2
XFILLER_194_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _05340_ _05341_ _04912_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__mux2_1
XFILLER_190_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _04351_ vssd1 vssd1 vccd1 vccd1 _04353_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19750_ rbzero.pov.spi_buffer\[14\] rbzero.pov.spi_buffer\[15\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16962_ _09981_ _09983_ vssd1 vssd1 vccd1 vccd1 _09984_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12085_ gpout0.vpos\[4\] _04418_ _04578_ _04652_ _05273_ vssd1 vssd1 vccd1 vccd1
+ _05274_ sky130_fd_sc_hd__a221o_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18701_ _02897_ _02898_ _02899_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21o_1
X_15913_ _08335_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__clkbuf_4
X_11036_ rbzero.tex_b1\[19\] rbzero.tex_b1\[20\] _04314_ vssd1 vssd1 vccd1 vccd1 _04317_
+ sky130_fd_sc_hd__mux2_1
X_16893_ _09913_ _09914_ vssd1 vssd1 vccd1 vccd1 _09915_ sky130_fd_sc_hd__nand2_1
XFILLER_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15844_ _08916_ _08937_ _08938_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__a21boi_1
X_18632_ _05127_ rbzero.wall_tracer.rayAddendY\[2\] _02813_ vssd1 vssd1 vccd1 vccd1
+ _02836_ sky130_fd_sc_hd__o21bai_1
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15775_ _08839_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__xor2_1
X_18563_ rbzero.debug_overlay.vplaneY\[-7\] _02764_ vssd1 vssd1 vccd1 vccd1 _02773_
+ sky130_fd_sc_hd__or2_1
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12987_ rbzero.wall_tracer.trackDistY\[9\] _06162_ vssd1 vssd1 vccd1 vccd1 _06163_
+ sky130_fd_sc_hd__or2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _01724_ _01719_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__or2b_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07872_ _07858_ _07827_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__mux2_1
X_11938_ rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__buf_2
X_18494_ rbzero.map_rom.a6 _02714_ _02704_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _01715_ _01737_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14657_ _06758_ _07331_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__and2_1
XFILLER_127_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11869_ reg_rgb\[6\] _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__mux2_2
XFILLER_159_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13608_ _06774_ _06777_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__and3_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17376_ _10150_ _10275_ _10280_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14588_ _07423_ _07444_ _07754_ _07758_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__o31a_1
X_16327_ _09417_ _09418_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__xnor2_1
X_19115_ _03110_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__clkbuf_4
X_13539_ _06709_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19046_ _05270_ _03091_ _03093_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__nand3_4
XFILLER_118_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _09238_ _09232_ _09349_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__and3_1
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15209_ _08164_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16189_ _08368_ _08814_ _09151_ _09281_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__o31a_1
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19948_ rbzero.debug_overlay.playerX\[4\] _03598_ vssd1 vssd1 vccd1 vccd1 _03604_
+ sky130_fd_sc_hd__nor2_1
XFILLER_136_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19879_ rbzero.pov.ss_buffer\[1\] rbzero.pov.ss_buffer\[0\] _03084_ vssd1 vssd1 vccd1
+ vccd1 _03552_ sky130_fd_sc_hd__mux2_1
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21910_ net436 _01499_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21841_ net367 _01430_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21772_ net298 _01361_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20723_ _03728_ clknet_1_0__leaf__05761_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__and2_2
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20654_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20585_ _09732_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__buf_4
XFILLER_176_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21206_ clknet_leaf_11_i_clk _00795_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21137_ clknet_leaf_31_i_clk _00726_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21068_ clknet_leaf_83_i_clk _00657_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20019_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__buf_2
X_12910_ rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__inv_2
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _06851_ _06875_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__and2b_1
XFILLER_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20503__348 clknet_1_0__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__inv_2
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12841_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _06013_
+ _06016_ _06011_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a221o_1
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _08172_ _08366_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__nand2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__inv_2
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _07676_ _07679_ _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _04892_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__buf_6
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _08585_ _08507_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__xnor2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17230_ _10017_ _10003_ _10121_ vssd1 vssd1 vccd1 vccd1 _10250_ sky130_fd_sc_hd__a21o_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _07608_ _07612_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__xor2_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11654_ rbzero.row_render.size\[7\] _04840_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _04090_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__clkbuf_1
X_17161_ _10081_ _10085_ vssd1 vssd1 vccd1 vccd1 _10181_ sky130_fd_sc_hd__and2b_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14373_ _07316_ _07443_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__or2_1
X_11585_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _04775_ sky130_fd_sc_hd__or2_1
XFILLER_128_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ _09203_ _09205_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13324_ _06370_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__inv_2
X_17092_ _09992_ _10024_ _10112_ vssd1 vssd1 vccd1 vccd1 _10113_ sky130_fd_sc_hd__a21oi_1
X_10536_ _03971_ _04051_ _04052_ _03977_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__or4b_4
XFILLER_182_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _09081_ _09075_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__and2b_1
XFILLER_115_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _06284_ _06320_ _06321_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__o21a_1
XFILLER_109_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10467_ rbzero.tex_r1\[31\] rbzero.tex_r1\[32\] _04013_ vssd1 vssd1 vccd1 vccd1 _04016_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ rbzero.tex_g1\[7\] _05305_ _05392_ _04947_ vssd1 vssd1 vccd1 vccd1 _05393_
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _06305_ _06307_ _06293_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__a21o_1
X_10398_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__buf_4
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19802_ _03467_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__buf_4
X_12137_ rbzero.tex_g0\[26\] _04924_ _04982_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a21o_1
XFILLER_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17994_ _01922_ _09195_ _02191_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o31a_1
XFILLER_150_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19733_ net511 rbzero.pov.spi_buffer\[7\] _03468_ vssd1 vssd1 vccd1 vccd1 _03476_
+ sky130_fd_sc_hd__mux2_1
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16945_ _09681_ _09966_ vssd1 vssd1 vccd1 vccd1 _09967_ sky130_fd_sc_hd__xnor2_2
X_12068_ rbzero.tex_r1\[50\] _05031_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__or2_1
XFILLER_81_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11019_ rbzero.tex_b1\[27\] rbzero.tex_b1\[28\] _04303_ vssd1 vssd1 vccd1 vccd1 _04308_
+ sky130_fd_sc_hd__mux2_1
X_16876_ _09659_ _09645_ vssd1 vssd1 vccd1 vccd1 _09898_ sky130_fd_sc_hd__or2b_1
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18615_ _09753_ _02812_ _02813_ _02820_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__a31o_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _08039_ _08274_ _08296_ _08458_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__or4_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ _03426_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15758_ _08852_ _08850_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__xnor2_1
X_18546_ rbzero.wall_tracer.rayAddendY\[-5\] _02606_ _09753_ _02755_ _02757_ vssd1
+ vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a221o_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14709_ _06613_ _07805_ _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15689_ _08743_ _08745_ _08744_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__a21o_1
XFILLER_127_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18477_ rbzero.wall_tracer.rayAddendX\[10\] _02701_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02702_ sky130_fd_sc_hd__mux2_1
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _08889_ _10330_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XFILLER_186_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17359_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _10377_ sky130_fd_sc_hd__nand2_1
XFILLER_140_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19029_ rbzero.map_overlay.i_otherx\[3\] _03101_ vssd1 vssd1 vccd1 vccd1 _03106_
+ sky130_fd_sc_hd__or2_1
X_22040_ clknet_leaf_37_i_clk _01629_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21824_ net350 _01413_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21755_ net281 _01344_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20706_ _03919_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nor2_1
XFILLER_197_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21686_ clknet_leaf_3_i_clk _01275_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20637_ _03861_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__xor2_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11370_ rbzero.spi_registers.texadd0\[22\] _04535_ _04561_ vssd1 vssd1 vccd1 vccd1
+ _04562_ sky130_fd_sc_hd__o21ai_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _06164_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 _06216_
+ sky130_fd_sc_hd__and2_1
XFILLER_156_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14991_ _08105_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13942_ _07072_ _07071_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__or2b_1
X_16730_ _06113_ _09118_ _09767_ vssd1 vssd1 vccd1 vccd1 _09768_ sky130_fd_sc_hd__a21o_1
XFILLER_207_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16661_ _09741_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__clkbuf_1
X_13873_ _07023_ _07029_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ _08695_ _08705_ _08706_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__a21oi_1
X_18400_ _02629_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__and2_1
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12824_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__and2_1
X_16592_ _08431_ _09559_ _09680_ _08733_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__a2bb2o_1
X_19380_ _02481_ rbzero.spi_registers.new_sky\[1\] _03309_ vssd1 vssd1 vccd1 vccd1
+ _03311_ sky130_fd_sc_hd__mux2_1
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _08404_ _08472_ _08637_ _08380_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__a2bb2o_1
X_18331_ rbzero.wall_tracer.rayAddendX\[-1\] _09745_ _02566_ _02534_ vssd1 vssd1 vccd1
+ vccd1 _02567_ sky130_fd_sc_hd__a22o_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12755_ _05888_ _05881_ _05053_ _05909_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__and4_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11706_ rbzero.floor_leak\[3\] _04889_ _04890_ rbzero.floor_leak\[2\] _04895_ vssd1
+ vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__o221a_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ rbzero.spi_registers.new_texadd\[2\]\[20\] rbzero.spi_registers.spi_buffer\[20\]
+ _02478_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15474_ _08547_ _08548_ _08567_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__nand3_1
XFILLER_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12686_ _04589_ _04704_ _04419_ _03973_ _05822_ net23 vssd1 vssd1 vccd1 vccd1 _05865_
+ sky130_fd_sc_hd__mux4_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17213_ _10231_ _10232_ vssd1 vssd1 vccd1 vccd1 _10233_ sky130_fd_sc_hd__nor2_1
XFILLER_129_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14425_ _07206_ _07476_ _07444_ _06720_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__o22a_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11637_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__buf_4
X_18193_ _02457_ _02458_ _06104_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a21o_1
XFILLER_156_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17144_ _09520_ _09252_ vssd1 vssd1 vccd1 vccd1 _10164_ sky130_fd_sc_hd__nor2_1
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14356_ _07472_ _07526_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__03782_ clknet_0__03782_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03782_
+ sky130_fd_sc_hd__clkbuf_16
X_11568_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _04758_ sky130_fd_sc_hd__or2_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ _06350_ _06352_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__nand2_2
X_10519_ rbzero.tex_r1\[6\] rbzero.tex_r1\[7\] _04035_ vssd1 vssd1 vccd1 vccd1 _04043_
+ sky130_fd_sc_hd__mux2_1
X_17075_ _10095_ vssd1 vssd1 vccd1 vccd1 _10096_ sky130_fd_sc_hd__buf_2
XFILLER_157_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14287_ _07452_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__xnor2_1
X_11499_ gpout0.vpos\[0\] _04686_ rbzero.debug_overlay.playerX\[-1\] _04446_ _04688_
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o221a_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _09120_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__buf_2
X_13238_ _06393_ _06406_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__and3_1
XFILLER_170_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13169_ _06319_ _06318_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__and2b_1
XFILLER_112_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17977_ _02263_ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__nor2_1
XFILLER_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19716_ _03440_ _03439_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__nand2_1
X_16928_ _09946_ _09948_ vssd1 vssd1 vccd1 vccd1 _09950_ sky130_fd_sc_hd__nand2_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16859_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09882_ sky130_fd_sc_hd__and2_1
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19578_ _03417_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18529_ rbzero.wall_tracer.mapX\[5\] _02741_ _09844_ vssd1 vssd1 vccd1 vccd1 _02742_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21540_ clknet_leaf_71_i_clk _01129_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ net189 _01060_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22023_ clknet_leaf_55_i_clk _01612_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _04226_ vssd1 vssd1 vccd1 vccd1 _04230_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21807_ net333 _01396_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ net13 net12 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__nor2_1
X_21738_ net264 _01327_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__buf_2
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21669_ clknet_leaf_32_i_clk _01258_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14210_ _07253_ _07331_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__nor2_1
XFILLER_32_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11422_ rbzero.spi_registers.texadd2\[1\] _04537_ _04457_ rbzero.spi_registers.texadd3\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a22o_1
XFILLER_177_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15190_ rbzero.wall_tracer.visualWallDist\[-3\] _08161_ vssd1 vssd1 vccd1 vccd1 _08285_
+ sky130_fd_sc_hd__or2_1
XFILLER_126_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14141_ _07308_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__xor2_1
X_11353_ _04461_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _07216_ _07217_ _07241_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nor3_1
XFILLER_180_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11284_ rbzero.spi_registers.texadd0\[11\] _04467_ _04474_ _04475_ vssd1 vssd1 vccd1
+ vccd1 _04476_ sky130_fd_sc_hd__o22a_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17900_ _02033_ _02092_ _02098_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__o21a_1
XFILLER_117_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13023_ rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__inv_2
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18880_ rbzero.pov.spi_buffer\[48\] rbzero.pov.ready_buffer\[48\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17831_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__xor2_1
X_20509__354 clknet_1_1__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__inv_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17762_ _01928_ _02050_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__o21ba_1
XFILLER_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14974_ _08096_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19501_ _03377_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
X_20360__219 clknet_1_1__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__inv_2
X_16713_ rbzero.traced_texa\[5\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__a22o_1
X_13925_ _07094_ _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_1
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17693_ _01983_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19432_ _02483_ rbzero.spi_registers.new_other\[2\] _03338_ vssd1 vssd1 vccd1 vccd1
+ _03341_ sky130_fd_sc_hd__mux2_1
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13856_ _06737_ _06808_ _06974_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__a21oi_1
X_16644_ _09731_ vssd1 vssd1 vccd1 vccd1 _09732_ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _05711_ _05952_ _05948_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__and3_1
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19363_ rbzero.spi_registers.new_vshift\[1\] _03297_ _03300_ _03278_ vssd1 vssd1
+ vccd1 vccd1 _00898_ sky130_fd_sc_hd__o211a_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16575_ _09167_ _09186_ _09556_ vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__or3_1
X_13787_ _06911_ _06956_ _06955_ _06946_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__o211a_1
X_10999_ _04297_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18314_ _02547_ _02548_ _02550_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__or3_1
X_15526_ _08616_ _08538_ _08620_ _08539_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__o31a_1
X_12738_ _05901_ _05908_ _05909_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a211o_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ rbzero.spi_registers.new_texadd\[3\]\[14\] _03254_ _03260_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__o211a_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15457_ _08304_ _08541_ _08551_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__or3_1
XFILLER_148_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18245_ _02497_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__clkbuf_1
X_12669_ _05053_ _05846_ _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__and3_1
XFILLER_124_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14408_ _07577_ _07578_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__and2_1
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20254__124 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__inv_2
X_15388_ _08481_ _08482_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18176_ _02443_ _02444_ _01981_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a21bo_1
XFILLER_11_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17127_ _10040_ _10053_ _10051_ vssd1 vssd1 vccd1 vccd1 _10147_ sky130_fd_sc_hd__a21o_1
X_14339_ _07424_ _07506_ _07509_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17058_ _08431_ _09560_ vssd1 vssd1 vccd1 vccd1 _10079_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__03796_ _03796_ vssd1 vssd1 vccd1 vccd1 clknet_0__03796_ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _09101_ _09103_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20971_ clknet_leaf_59_i_clk _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21523_ clknet_leaf_84_i_clk _01112_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21454_ net172 _01043_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21385_ clknet_leaf_23_i_clk _00974_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19694__72 clknet_1_0__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
XFILLER_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__buf_2
XFILLER_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22006_ net128 _01595_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20198_ rbzero.spi_registers.new_texadd\[3\]\[14\] rbzero.spi_registers.spi_buffer\[14\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__mux2_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11971_ rbzero.debug_overlay.playerX\[5\] _05101_ _05112_ rbzero.debug_overlay.playerX\[-5\]
+ _04646_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a221o_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03785_ clknet_0__03785_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03785_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _06878_ _06880_ _06774_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__a21boi_1
X_10922_ rbzero.tex_g0\[10\] rbzero.tex_g0\[9\] _04248_ vssd1 vssd1 vccd1 vccd1 _04257_
+ sky130_fd_sc_hd__mux2_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _07827_ _07858_ _07860_ _07822_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__a211o_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13641_ _06804_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__xor2_1
X_10853_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _04215_ vssd1 vssd1 vccd1 vccd1 _04221_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _09405_ _09451_ vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__xnor2_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _06682_ _06737_ _06728_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__a21o_1
XFILLER_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10784_ _04184_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15311_ rbzero.wall_tracer.stepDistY\[-1\] _08405_ vssd1 vssd1 vccd1 vccd1 _08406_
+ sky130_fd_sc_hd__nand2_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ net10 vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__buf_2
X_16291_ _09361_ _09382_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15242_ _08336_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__clkbuf_4
X_18030_ _02309_ _02316_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__xnor2_1
X_12454_ _05636_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _04489_ _04499_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__xnor2_1
X_15173_ _08266_ _08267_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__nand2_1
XFILLER_158_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _05009_ vssd1 vssd1 vccd1 vccd1 _05570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _07293_ _07294_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11336_ rbzero.spi_registers.texadd1\[16\] _04461_ _04470_ _04527_ vssd1 vssd1 vccd1
+ vccd1 _04528_ sky130_fd_sc_hd__a211o_1
XFILLER_181_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19981_ _08309_ _03561_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nor2_1
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18932_ rbzero.pov.spi_buffer\[73\] rbzero.pov.ready_buffer\[73\] _02967_ vssd1 vssd1
+ vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
X_14055_ _06640_ _06769_ _07185_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__nor3_1
X_11267_ rbzero.wall_hot\[1\] vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__inv_2
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13006_ rbzero.wall_tracer.trackDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__inv_2
X_18863_ _03012_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11198_ _04401_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17814_ _01922_ _09315_ _02101_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18794_ rbzero.pov.spi_buffer\[7\] rbzero.pov.ready_buffer\[7\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
X_17745_ _01832_ _02030_ _02033_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__nand3_1
XFILLER_130_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14957_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.trackDistX\[8\] _06217_
+ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__mux2_1
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13908_ _06748_ _06721_ _07078_ _06732_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__o2bb2a_1
X_17676_ _01965_ _01966_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and2_1
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14888_ _06217_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__buf_4
XFILLER_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19415_ _03331_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ _09714_ _09716_ vssd1 vssd1 vccd1 vccd1 _09717_ sky130_fd_sc_hd__nor2_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13839_ _06926_ _06970_ _06966_ _06969_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a211o_1
XFILLER_189_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ rbzero.color_floor\[0\] _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
X_16558_ _08535_ _08409_ _09647_ _08152_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__o22ai_1
XFILLER_204_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _08172_ _08305_ _08352_ _08350_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__a31o_1
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19277_ rbzero.spi_registers.new_texadd\[3\]\[7\] _03240_ _03250_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00862_ sky130_fd_sc_hd__o211a_1
X_16489_ _09578_ _09579_ vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__nor2_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18228_ rbzero.spi_registers.new_texadd\[2\]\[4\] _02487_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18159_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__or2_1
XFILLER_190_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21170_ clknet_leaf_14_i_clk _00759_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20121_ _03715_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__03779_ _03779_ vssd1 vssd1 vccd1 vccd1 clknet_0__03779_ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20052_ rbzero.debug_overlay.facingY\[-7\] _03676_ _03677_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01210_ sky130_fd_sc_hd__a211o_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ clknet_leaf_65_i_clk _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ clknet_leaf_44_i_clk _00474_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20538__380 clknet_1_1__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__inv_2
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21506_ clknet_leaf_98_i_clk _01095_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21437_ net155 _01026_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12170_ rbzero.tex_g0\[50\] _04924_ _04982_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a21o_1
X_21368_ clknet_leaf_12_i_clk _00957_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _04351_ vssd1 vssd1 vccd1 vccd1 _04361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21299_ clknet_leaf_30_i_clk _00888_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _03978_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _08952_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__o21ba_1
XFILLER_153_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20283__150 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__inv_2
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14811_ _06619_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__and3_1
XFILLER_188_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _08873_ _08878_ _08885_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__o21ai_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _01818_ _09186_ _01706_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o31a_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ rbzero.debug_overlay.facingY\[10\] _05105_ _05142_ vssd1 vssd1 vccd1 vccd1
+ _05143_ sky130_fd_sc_hd__a21oi_2
X_14742_ _07827_ _07805_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__and2_1
Xtop_ew_algofoogle_104 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_104/HI zeros[11]
+ sky130_fd_sc_hd__conb_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_115 vssd1 vssd1 vccd1 vccd1 ones[6] top_ew_algofoogle_115/LO sky130_fd_sc_hd__conb_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _04214_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__clkbuf_4
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17461_ _01752_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__xor2_4
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14673_ _07402_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__clkinv_2
XFILLER_189_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11885_ _04421_ _04636_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__nor2_1
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19200_ rbzero.spi_registers.got_new_texadd\[2\] _03096_ vssd1 vssd1 vccd1 vccd1
+ _03205_ sky130_fd_sc_hd__nand2_2
X_16412_ _09388_ _09390_ _09502_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__a21oi_1
X_13624_ _06791_ _06793_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__or2_1
X_10836_ _04211_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ _01683_ _01684_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nor2_1
XFILLER_73_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19131_ rbzero.spi_registers.texadd0\[18\] _03156_ vssd1 vssd1 vccd1 vccd1 _03166_
+ sky130_fd_sc_hd__or2_1
XFILLER_201_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16343_ _09307_ _09312_ _09434_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__a21bo_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ _06692_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__buf_4
X_10767_ _04175_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ clknet_3_3_0_i_clk _05664_ _05638_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__and3_2
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16274_ _08616_ _09363_ _09365_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__o21ba_1
XFILLER_121_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19062_ rbzero.map_overlay.i_mapdx\[4\] _03122_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__or2_1
XFILLER_158_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _06594_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__and2_2
XFILLER_157_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ rbzero.tex_g1\[51\] rbzero.tex_g1\[52\] _04132_ vssd1 vssd1 vccd1 vccd1 _04139_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18013_ _01922_ _09433_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__nor2_1
X_15225_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerY\[-2\] _08281_
+ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__or3_2
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ _04817_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__or2_1
XFILLER_201_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15156_ rbzero.wall_tracer.stepDistX\[-6\] _06261_ vssd1 vssd1 vccd1 vccd1 _08251_
+ sky130_fd_sc_hd__or2_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12368_ rbzero.color_sky\[5\] rbzero.color_floor\[5\] _04825_ vssd1 vssd1 vccd1 vccd1
+ _05553_ sky130_fd_sc_hd__mux2_1
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14107_ _07187_ _07231_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__a21bo_1
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11319_ _04464_ _04472_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__nor2_1
XFILLER_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19964_ net41 _03557_ _03095_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__o21a_1
X_15087_ _06402_ _06349_ _08181_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__and3_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19673__53 clknet_1_1__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
X_12299_ rbzero.tex_b0\[55\] _04926_ _04928_ _04891_ vssd1 vssd1 vccd1 vccd1 _05485_
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14038_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__clkbuf_4
X_18915_ _03039_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
X_20366__225 clknet_1_1__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__inv_2
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03464_ clknet_0__03464_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03464_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19895_ _03559_ _03562_ _03563_ _03302_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__o211a_1
XFILLER_68_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18846_ _03003_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18777_ rbzero.pov.spi_done _08116_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_209_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15989_ _08622_ _09082_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__or2_1
XFILLER_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17728_ _02016_ _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nor2_1
XFILLER_208_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _01842_ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20670_ _03888_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21o_1
XFILLER_189_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19329_ rbzero.spi_registers.got_new_sky _03097_ vssd1 vssd1 vccd1 vccd1 _03280_
+ sky130_fd_sc_hd__nand2_2
XFILLER_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21222_ clknet_leaf_28_i_clk _00811_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21153_ clknet_leaf_4_i_clk _00742_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20104_ _05129_ _03655_ _03706_ _03695_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__a211o_1
XFILLER_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21084_ clknet_leaf_88_i_clk _00673_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20035_ rbzero.pov.ready_buffer\[39\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03668_
+ sky130_fd_sc_hd__and3_1
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21986_ net132 _01575_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ clknet_leaf_48_i_clk _00526_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11670_ gpout0.hpos\[4\] _04850_ _04849_ _04411_ _04859_ vssd1 vssd1 vccd1 vccd1
+ _04860_ sky130_fd_sc_hd__o221a_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ clknet_leaf_20_i_clk _00457_ vssd1 vssd1 vccd1 vccd1 reg_rgb\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10621_ _04098_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20799_ clknet_leaf_47_i_clk _00388_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ _06379_ _06414_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__nand2_1
X_10552_ _04062_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _06421_ _06438_ _06441_ _06415_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__o211ai_1
X_10483_ _03979_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ rbzero.wall_tracer.stepDistX\[10\] _08031_ _08091_ vssd1 vssd1 vccd1 vccd1
+ _08115_ sky130_fd_sc_hd__mux2_1
X_12222_ rbzero.tex_g1\[16\] _05185_ _05181_ _05407_ _05408_ vssd1 vssd1 vccd1 vccd1
+ _05409_ sky130_fd_sc_hd__a311o_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20315__179 clknet_1_0__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__inv_2
XFILLER_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _04948_ vssd1 vssd1 vccd1 vccd1 _05341_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _04352_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16961_ _09684_ _09696_ _09982_ vssd1 vssd1 vccd1 vccd1 _09983_ sky130_fd_sc_hd__a21o_1
X_12084_ _04648_ _04411_ _04578_ _04652_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__o22ai_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18700_ _02897_ _02898_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__nand3_1
X_15912_ _09004_ _09006_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__nand2_1
X_11035_ _04316_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16892_ _08731_ _09079_ _09628_ vssd1 vssd1 vccd1 vccd1 _09914_ sky130_fd_sc_hd__or3_1
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ rbzero.wall_tracer.rayAddendY\[2\] rbzero.wall_tracer.rayAddendY\[1\] _05127_
+ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o21ai_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _08917_ _08936_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__or2_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _02767_ _02768_ _02770_ _02771_ _04442_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__o311a_1
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _08856_ _08855_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__or2b_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12986_ rbzero.wall_tracer.trackDistX\[9\] vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__inv_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _01708_ _01709_ _01711_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__o21ai_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _06589_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__buf_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ rbzero.debug_overlay.vplaneX\[10\] _05105_ _05109_ _05125_ vssd1 vssd1 vccd1
+ vccd1 _05126_ sky130_fd_sc_hd__a211o_2
X_18493_ rbzero.debug_overlay.playerY\[3\] _02713_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02714_ sky130_fd_sc_hd__mux2_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _01734_ _01736_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__xor2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11868_ net45 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__buf_6
X_14656_ _06613_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__buf_2
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10819_ _04202_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13607_ _06681_ _06775_ _06776_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a21o_1
X_17375_ _01666_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__nand2_1
X_11799_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _04948_ vssd1 vssd1 vccd1 vccd1 _04989_
+ sky130_fd_sc_hd__mux2_1
X_14587_ _07755_ _07757_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nand2_1
XFILLER_203_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19114_ rbzero.spi_registers.texadd0\[10\] _03156_ vssd1 vssd1 vccd1 vccd1 _03157_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16326_ _09315_ _09306_ _08431_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13538_ _06617_ _06640_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__or3b_1
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19045_ rbzero.spi_registers.got_new_vinf vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__inv_2
XFILLER_12_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13469_ _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__buf_4
X_16257_ _09238_ _09232_ _09349_ vssd1 vssd1 vccd1 vccd1 _09350_ sky130_fd_sc_hd__a21oi_1
XFILLER_199_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15208_ _08238_ _08289_ _08302_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__a21bo_1
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04634_ clknet_0__04634_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04634_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16188_ _09153_ _09154_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__nand2_1
XFILLER_160_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15139_ _08229_ _08233_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__or2_1
XFILLER_5_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19947_ _03559_ _03599_ rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1
+ _03603_ sky130_fd_sc_hd__o21a_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19878_ _03551_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18829_ _02994_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21840_ net366 _01429_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21771_ net297 _01360_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20420__274 clknet_1_0__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__inv_2
X_20722_ _03931_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__buf_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20653_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03876_
+ sky130_fd_sc_hd__or2_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20584_ _03734_ _03817_ _03818_ _03814_ rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1
+ _01601_ sky130_fd_sc_hd__a32o_1
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21205_ clknet_leaf_11_i_clk _00794_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21136_ clknet_leaf_32_i_clk _00725_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19652__34 clknet_1_0__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21067_ clknet_leaf_83_i_clk _00656_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20018_ _03095_ _03557_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__and2_1
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _06014_
+ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a31o_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20565__25 clknet_1_0__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ net36 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__buf_2
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ net495 _01558_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _04827_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__buf_4
X_14510_ _07647_ _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__or2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _08178_ _08213_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__nor2_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20395__251 clknet_1_1__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__inv_2
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14441_ _07609_ _07610_ _07611_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__a21boi_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__nor2_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _04088_ vssd1 vssd1 vccd1 vccd1 _04090_
+ sky130_fd_sc_hd__mux2_1
X_17160_ _10064_ _10072_ _10071_ vssd1 vssd1 vccd1 vccd1 _10180_ sky130_fd_sc_hd__a21o_1
XFILLER_161_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14372_ _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__inv_2
XFILLER_70_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19715__90 clknet_1_0__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
X_11584_ _04770_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _09041_ _09059_ _09204_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__a21bo_1
X_13323_ _06485_ _06491_ _06493_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__or3_2
XFILLER_156_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10535_ _03974_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__clkinv_4
X_17091_ _10056_ _10111_ vssd1 vssd1 vccd1 vccd1 _10112_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16042_ _09134_ _09135_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__nand2_1
XFILLER_170_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13254_ _06416_ _06417_ _06418_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__or4b_1
X_10466_ _04015_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ rbzero.tex_g1\[6\] _04831_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or2_1
XFILLER_142_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _04443_ _06353_ _06354_ _06355_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__o2bb2a_4
X_10397_ _03971_ _03973_ _03974_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and4_2
X_19801_ _03511_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
X_12136_ rbzero.tex_g0\[27\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__and3_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ _02189_ _02190_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__nand2_1
X_19732_ _03475_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
X_16944_ _08910_ _09559_ vssd1 vssd1 vccd1 vccd1 _09966_ sky130_fd_sc_hd__nor2_1
X_12067_ rbzero.tex_r1\[52\] _05199_ _04924_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _04307_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16875_ _09623_ _09636_ _09635_ vssd1 vssd1 vccd1 vccd1 _09897_ sky130_fd_sc_hd__a21o_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18614_ rbzero.wall_tracer.rayAddendY\[1\] _09744_ _02819_ _02534_ vssd1 vssd1 vccd1
+ vccd1 _02820_ sky130_fd_sc_hd__a22o_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _08337_ _08441_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__nor2_1
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19594_ rbzero.spi_registers.new_texadd\[1\]\[14\] rbzero.spi_registers.spi_buffer\[14\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20478__326 clknet_1_1__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__inv_2
X_18545_ _02756_ _04442_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__nor2_1
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757_ _08843_ _08845_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__nand2_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ rbzero.map_overlay.i_mapdx\[0\] _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and2_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _06613_ _07809_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__nor2_1
X_18476_ _04434_ _02699_ _02700_ _02694_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a22o_1
X_15688_ _08748_ _08750_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__xnor2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _08816_ _10215_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__or2_1
XFILLER_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ _06579_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__nor2_1
XFILLER_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17358_ _06171_ _09785_ _10376_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _09396_ _09399_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__and2_1
XFILLER_174_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17289_ _10272_ _10307_ vssd1 vssd1 vccd1 vccd1 _10308_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19028_ rbzero.spi_registers.new_other\[8\] _03098_ _03105_ _03103_ vssd1 vssd1 vccd1
+ vccd1 _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21823_ net349 _01412_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21754_ net280 _01343_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20705_ _03914_ _03917_ _03918_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a21oi_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21685_ clknet_leaf_3_i_clk _01274_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20636_ _03854_ _03856_ _03855_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21boi_1
XFILLER_177_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21119_ clknet_leaf_70_i_clk _00708_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_14990_ rbzero.wall_tracer.stepDistX\[0\] _07992_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08105_ sky130_fd_sc_hd__mux2_1
XFILLER_93_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13941_ _07086_ _07098_ _07111_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16660_ _09739_ _09740_ _09732_ vssd1 vssd1 vccd1 vccd1 _09741_ sky130_fd_sc_hd__and3b_1
XFILLER_207_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13872_ _07011_ _07012_ _07014_ _07042_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a22o_1
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15611_ _08662_ _08694_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__nor2_1
X_12823_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__xnor2_1
X_16591_ _08431_ _09680_ vssd1 vssd1 vccd1 vccd1 _09681_ sky130_fd_sc_hd__nand2b_2
X_18330_ _05111_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__xor2_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15542_ _08581_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__inv_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _05884_ _05889_ _05931_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__and3_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ rbzero.floor_leak\[2\] _04814_ _04891_ rbzero.floor_leak\[1\] _04894_ vssd1
+ vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a221o_1
X_18261_ _02505_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__clkbuf_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15473_ _08547_ _08548_ _08567_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__a21o_1
X_12685_ net27 _05832_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__and3_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _10228_ _10230_ vssd1 vssd1 vccd1 vccd1 _10232_ sky130_fd_sc_hd__and2_1
X_11636_ _04786_ _04806_ _04815_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__nor3b_4
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14424_ _07590_ _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__or2_1
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18192_ _02457_ _02458_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__nor2_1
XFILLER_129_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17143_ _10161_ _10162_ vssd1 vssd1 vccd1 vccd1 _10163_ sky130_fd_sc_hd__nand2_1
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _04757_ sky130_fd_sc_hd__nand2_1
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14355_ _07524_ _07525_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__03781_ clknet_0__03781_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03781_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ _04042_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13306_ _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__xnor2_2
X_17074_ _08950_ _08581_ _09691_ _10093_ _10094_ vssd1 vssd1 vccd1 vccd1 _10095_ sky130_fd_sc_hd__o41a_1
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14286_ _07455_ _07456_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__xor2_1
X_11498_ _04687_ rbzero.debug_overlay.playerY\[-1\] vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _06087_ _09119_ _08395_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__mux2_1
X_13237_ _06324_ _06328_ _06407_ _06322_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__a31oi_4
X_10449_ _04006_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13168_ _06285_ _06287_ _06317_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__and3_1
XFILLER_112_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12119_ rbzero.tex_g0\[3\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__and3_1
X_13099_ rbzero.map_rom.i_row\[4\] rbzero.wall_tracer.mapY\[5\] rbzero.wall_tracer.mapY\[7\]
+ rbzero.wall_tracer.mapY\[6\] _06077_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__o41a_1
X_17976_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__nor2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16927_ _09946_ _09948_ vssd1 vssd1 vccd1 vccd1 _09949_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_62_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09881_ sky130_fd_sc_hd__nor2_1
XFILLER_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15809_ _08864_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__nor2_1
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19577_ rbzero.spi_registers.new_texadd\[1\]\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__mux2_1
XFILLER_207_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16789_ _09817_ _09818_ _09819_ vssd1 vssd1 vccd1 vccd1 _09820_ sky130_fd_sc_hd__and3_1
XFILLER_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_77_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_197_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18528_ rbzero.debug_overlay.playerX\[5\] _02740_ _08123_ vssd1 vssd1 vccd1 vccd1
+ _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18459_ _02673_ _02674_ _02684_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__nand3_1
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21470_ net188 _01059_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20532__375 clknet_1_0__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__inv_2
XFILLER_147_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20231__103 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__inv_2
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22022_ clknet_leaf_54_i_clk _01611_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21806_ net332 _01395_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21737_ net263 _01326_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12470_ gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__clkbuf_4
XFILLER_138_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21668_ clknet_leaf_32_i_clk _01257_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _04575_ _04612_ _04452_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20619_ _03844_ _03845_ _03846_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a21o_1
X_21599_ clknet_leaf_70_i_clk _01188_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14140_ _06758_ _07310_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__and2_1
XFILLER_125_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _04534_ _04540_ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__and3_1
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14071_ _07216_ _07217_ _07241_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__o21a_2
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ rbzero.spi_registers.texadd3\[11\] _04465_ _04456_ rbzero.spi_registers.texadd2\[11\]
+ _04470_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a221o_1
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _06179_ rbzero.wall_tracer.trackDistX\[-2\] vssd1 vssd1 vccd1 vccd1 _06198_
+ sky130_fd_sc_hd__or2_1
XFILLER_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17830_ _02041_ _02060_ _02039_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17761_ _09528_ _10215_ _01718_ _08814_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__o22a_1
X_14973_ rbzero.wall_tracer.stepDistX\[-8\] _07923_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08096_ sky130_fd_sc_hd__mux2_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19500_ rbzero.spi_registers.new_mapd\[14\] rbzero.spi_registers.spi_buffer\[14\]
+ _03361_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__mux2_1
XFILLER_208_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ rbzero.traced_texa\[4\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a22o_1
XFILLER_130_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13924_ _06770_ _06877_ _07093_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__a21oi_1
X_17692_ rbzero.wall_tracer.trackDistX\[6\] _01982_ _09844_ vssd1 vssd1 vccd1 vccd1
+ _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19431_ _03340_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16643_ _04408_ _09729_ vssd1 vssd1 vccd1 vccd1 _09731_ sky130_fd_sc_hd__nor2_1
X_13855_ _06982_ _06681_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__nand2_1
X_12806_ net53 _05944_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a21o_1
X_19362_ rbzero.spi_registers.vshift\[1\] _03298_ vssd1 vssd1 vccd1 vccd1 _03300_
+ sky130_fd_sc_hd__or2_1
X_16574_ _09410_ _09663_ _09550_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__a21bo_1
X_10998_ rbzero.tex_b1\[37\] rbzero.tex_b1\[38\] _04292_ vssd1 vssd1 vccd1 vccd1 _04297_
+ sky130_fd_sc_hd__mux2_1
X_13786_ _06946_ _06955_ _06956_ _06911_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a211oi_2
XFILLER_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18313_ _02538_ _02541_ _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15525_ _08553_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__clkbuf_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12737_ net31 _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nor2_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ rbzero.spi_registers.texadd3\[14\] _03255_ vssd1 vssd1 vccd1 vccd1 _03260_
+ sky130_fd_sc_hd__or2_1
XFILLER_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ rbzero.spi_registers.new_texadd\[2\]\[11\] rbzero.spi_registers.spi_buffer\[11\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
X_15456_ _08549_ _08550_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__and2_1
XFILLER_31_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14407_ _07473_ _07523_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__xor2_2
XFILLER_175_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18175_ _02440_ _02441_ _02442_ _08123_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__o31a_1
X_11619_ _04806_ _04807_ _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or3b_1
X_15387_ _08434_ _08384_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__nor2_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ net21 _05773_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__and3_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17126_ _10144_ _10145_ vssd1 vssd1 vccd1 vccd1 _10146_ sky130_fd_sc_hd__nor2_1
XFILLER_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14338_ _07507_ _07508_ _07426_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _09671_ _10077_ _09958_ _09959_ vssd1 vssd1 vccd1 vccd1 _10078_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_144_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03795_ _03795_ vssd1 vssd1 vccd1 vccd1 clknet_0__03795_ sky130_fd_sc_hd__clkbuf_16
X_14269_ _07438_ _07439_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__and2_1
XFILLER_143_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ _08220_ _09102_ _08138_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__mux2_1
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _02132_ _02133_ _02129_ _02131_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__o2bb2a_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20970_ clknet_leaf_59_i_clk _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19629_ rbzero.pov.spi_counter\[2\] _03442_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__and2_1
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21522_ clknet_leaf_84_i_clk _01111_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21453_ net171 _01042_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21384_ clknet_leaf_23_i_clk _00973_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20335_ clknet_1_1__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__buf_1
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__clkbuf_1
X_22005_ net127 _01594_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20197_ _03765_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11970_ rbzero.debug_overlay.playerX\[-8\] _05117_ _05122_ rbzero.debug_overlay.playerX\[-9\]
+ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
XFILLER_99_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03784_ clknet_0__03784_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03784_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ _04256_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10852_ _04220_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__clkbuf_1
X_13640_ _06806_ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__nand2_1
XFILLER_204_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10783_ rbzero.tex_g1\[11\] rbzero.tex_g1\[12\] _04177_ vssd1 vssd1 vccd1 vccd1 _04184_
+ sky130_fd_sc_hd__mux2_1
X_13571_ _06682_ _06693_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__nand2_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _08168_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__buf_4
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ net12 vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__inv_2
X_16290_ _09367_ _09381_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__xor2_1
X_20238__109 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__inv_2
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _08332_ _08335_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__or2_1
XFILLER_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ reg_hsync _05635_ _05058_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__mux2_2
XFILLER_200_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11404_ _04501_ _04503_ _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a21oi_1
X_12384_ _05199_ _05566_ _05568_ _04952_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o211a_1
X_15172_ _08235_ _08246_ _08253_ _08265_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__o22ai_1
XFILLER_158_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ rbzero.spi_registers.texadd3\[16\] _04526_ _04456_ rbzero.spi_registers.texadd2\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a22o_1
X_14123_ _07227_ _07271_ _07273_ _07270_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__o211a_1
XFILLER_180_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19980_ rbzero.debug_overlay.playerY\[-3\] _03617_ _03627_ _03579_ vssd1 vssd1 vccd1
+ vccd1 _01188_ sky130_fd_sc_hd__o211a_1
XFILLER_181_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18931_ _03047_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
X_11266_ rbzero.spi_registers.texadd2\[14\] _04456_ _04457_ rbzero.spi_registers.texadd3\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a22o_1
X_14054_ _06733_ _06769_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__or2_1
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _06179_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.trackDistX\[-3\]
+ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a22o_1
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18862_ rbzero.pov.spi_buffer\[39\] rbzero.pov.ready_buffer\[39\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
X_11197_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _04395_ vssd1 vssd1 vccd1 vccd1 _04401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _01922_ _09315_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__or3_1
XFILLER_122_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18793_ _02975_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17744_ _01832_ _02030_ _02033_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a21o_1
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14956_ _08065_ _08083_ _08084_ _08085_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__o211a_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13907_ _06710_ _06724_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__and2_1
X_17675_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__nand2_1
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14887_ _08035_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19414_ _02481_ rbzero.spi_registers.new_leak\[1\] _03329_ vssd1 vssd1 vccd1 vccd1
+ _03331_ sky130_fd_sc_hd__mux2_1
X_16626_ _09483_ _09585_ _09715_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13838_ _07005_ _07007_ _06963_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__a211oi_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19345_ rbzero.spi_registers.got_new_floor _03096_ vssd1 vssd1 vccd1 vccd1 _03290_
+ sky130_fd_sc_hd__and2_1
X_16557_ _08382_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__clkbuf_4
XFILLER_149_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13769_ _06933_ _06934_ _06939_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15508_ _08601_ _08602_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__nor2_1
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19276_ rbzero.spi_registers.texadd3\[7\] _03242_ vssd1 vssd1 vccd1 vccd1 _03250_
+ sky130_fd_sc_hd__or2_1
X_16488_ _09405_ _09451_ _09449_ vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__a21oi_1
X_18227_ rbzero.spi_registers.spi_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__buf_4
X_15439_ _08532_ _08533_ vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18158_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__nand2_1
XFILLER_156_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17109_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] _10015_
+ vssd1 vssd1 vccd1 vccd1 _10130_ sky130_fd_sc_hd__a21o_1
XFILLER_190_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18089_ _02366_ _02367_ _02368_ _06104_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a31o_1
XFILLER_137_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20120_ _02968_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__and2_1
XFILLER_172_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03778_ _03778_ vssd1 vssd1 vccd1 vccd1 clknet_0__03778_ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20051_ rbzero.pov.ready_buffer\[24\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__and3_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20343__204 clknet_1_0__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__inv_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ clknet_leaf_61_i_clk _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ clknet_leaf_44_i_clk _00473_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_202_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21505_ clknet_leaf_98_i_clk _01094_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21436_ net154 _01025_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21367_ clknet_leaf_12_i_clk _00956_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _04360_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21298_ clknet_leaf_31_i_clk _00887_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11051_ _04324_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14810_ _07972_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__clkbuf_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _08879_ _08884_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__nand2_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14741_ _07806_ _07858_ _07876_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__a21oi_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ rbzero.debug_overlay.facingY\[0\] _05115_ _05137_ _05141_ vssd1 vssd1 vccd1
+ vccd1 _05142_ sky130_fd_sc_hd__a211o_1
Xtop_ew_algofoogle_105 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_105/HI zeros[12]
+ sky130_fd_sc_hd__conb_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_116 vssd1 vssd1 vccd1 vccd1 ones[7] top_ew_algofoogle_116/LO sky130_fd_sc_hd__conb_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _10363_ _10364_ _10366_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__o21a_1
X_10904_ _04247_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _06720_ _07829_ _07828_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__a21oi_1
X_11884_ _05066_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__xor2_2
XFILLER_199_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16411_ _09498_ _09501_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13623_ _06791_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__xor2_1
X_17391_ _10287_ _10298_ _10296_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a21oi_1
X_10835_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _04203_ vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19130_ rbzero.spi_registers.new_texadd\[0\]\[17\] _03155_ _03165_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__o211a_1
X_16342_ _08461_ _09192_ _09433_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__or3_1
XFILLER_38_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13554_ _06710_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__nand2_2
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10766_ rbzero.tex_g1\[19\] rbzero.tex_g1\[20\] _04166_ vssd1 vssd1 vccd1 vccd1 _04175_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20439__290 clknet_1_0__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__inv_2
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19061_ rbzero.spi_registers.new_mapd\[13\] _03120_ _03126_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00770_ sky130_fd_sc_hd__o211a_1
X_12505_ _05658_ _04052_ _05638_ _05643_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__o211a_1
X_16273_ _08304_ _09243_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10697_ _04138_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ _06370_ _06590_ _06645_ _06584_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__o211a_1
X_18012_ _02195_ _02199_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a21o_1
X_15224_ rbzero.debug_overlay.playerY\[-1\] _06087_ vssd1 vssd1 vccd1 vccd1 _08319_
+ sky130_fd_sc_hd__nor2_1
X_12436_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _04892_ vssd1 vssd1 vccd1 vccd1 _05621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15155_ rbzero.wall_tracer.stepDistY\[-6\] _08157_ _08247_ _08249_ vssd1 vssd1 vccd1
+ vccd1 _08250_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_201_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12367_ _05552_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_153_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _07224_ _07230_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or2b_1
XFILLER_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11318_ _04481_ _04507_ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a21o_1
X_12298_ rbzero.tex_b0\[54\] _05314_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__and2_1
XFILLER_141_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15086_ _06353_ _06358_ _08180_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__and3_1
X_19963_ _03611_ _03614_ _03615_ _03579_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__o211a_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14037_ _07161_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__nand2_1
X_18914_ rbzero.pov.spi_buffer\[64\] rbzero.pov.ready_buffer\[64\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
X_11249_ _03977_ _04417_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__nand2_2
Xclkbuf_1_1__f__03463_ clknet_0__03463_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03463_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19894_ _03560_ _03559_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__nand2_1
X_18845_ rbzero.pov.spi_buffer\[31\] rbzero.pov.ready_buffer\[31\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03003_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18776_ _02965_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
X_15988_ _08622_ _09082_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__nand2_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17727_ _02015_ _02014_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__and2b_1
X_14939_ rbzero.wall_tracer.visualWallDist\[2\] _08046_ vssd1 vssd1 vccd1 vccd1 _08074_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17658_ _01941_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__xor2_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ _09558_ _09571_ _09698_ vssd1 vssd1 vccd1 vccd1 _09699_ sky130_fd_sc_hd__a21o_1
XFILLER_189_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _01878_ _01879_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nor2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19328_ rbzero.spi_registers.new_leak\[5\] _03271_ _03279_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00884_ sky130_fd_sc_hd__o211a_1
XFILLER_188_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19259_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21221_ clknet_leaf_28_i_clk _00810_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21152_ clknet_leaf_3_i_clk _00741_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20103_ rbzero.pov.ready_buffer\[3\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03706_
+ sky130_fd_sc_hd__and3_1
XFILLER_160_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21083_ clknet_leaf_88_i_clk _00672_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20034_ rbzero.debug_overlay.facingX\[-4\] _03663_ _03667_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01202_ sky130_fd_sc_hd__a211o_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ net131 _01574_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ clknet_leaf_49_i_clk _00525_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20867_ clknet_leaf_65_i_clk _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _04088_ vssd1 vssd1 vccd1 vccd1 _04098_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20798_ clknet_leaf_47_i_clk _00387_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10551_ rbzero.tex_r0\[58\] rbzero.tex_r0\[57\] _04055_ vssd1 vssd1 vccd1 vccd1 _04062_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10482_ _04023_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__clkbuf_1
X_13270_ _06322_ _06419_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nor2_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ rbzero.tex_g1\[17\] _04905_ _05186_ _04919_ vssd1 vssd1 vccd1 vccd1 _05408_
+ sky130_fd_sc_hd__a31o_1
XFILLER_68_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21419_ clknet_leaf_4_i_clk _01008_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12152_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _05010_ vssd1 vssd1 vccd1 vccd1 _05340_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11103_ rbzero.tex_b0\[52\] rbzero.tex_b0\[51\] _04351_ vssd1 vssd1 vccd1 vccd1 _04352_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16960_ _09693_ _09695_ vssd1 vssd1 vccd1 vccd1 _09982_ sky130_fd_sc_hd__nor2_1
X_12083_ _04656_ _04628_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _08151_ _09005_ _08952_ _08166_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__o22ai_1
X_11034_ rbzero.tex_b1\[20\] rbzero.tex_b1\[21\] _04314_ vssd1 vssd1 vccd1 vccd1 _04316_
+ sky130_fd_sc_hd__mux2_1
X_16891_ _09525_ _09079_ _09628_ vssd1 vssd1 vccd1 vccd1 _09913_ sky130_fd_sc_hd__o21ai_1
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18630_ _05127_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02834_
+ sky130_fd_sc_hd__nor2_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _08917_ _08936_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__xor2_1
XFILLER_65_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _02767_ _02768_ _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o21ai_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _08830_ _08861_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__xor2_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ _06106_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__nand2_2
XFILLER_205_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17512_ _01772_ _01803_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__xnor2_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _07893_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__clkbuf_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ rbzero.debug_overlay.vplaneX\[-3\] _05110_ _05114_ _05124_ vssd1 vssd1 vccd1
+ vccd1 _05125_ sky130_fd_sc_hd__a211o_1
X_18492_ _06095_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__xnor2_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _10339_ _10347_ _01735_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14655_ _06595_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__buf_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ rbzero.trace_state\[0\] _04635_ _05052_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_
+ sky130_fd_sc_hd__o211a_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__05820_ clknet_0__05820_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05820_
+ sky130_fd_sc_hd__clkbuf_16
X_13606_ _06729_ _06775_ _06776_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__and3_1
X_17374_ _09525_ _09491_ _01665_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__o21ai_1
X_10818_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _04121_ vssd1 vssd1 vccd1 vccd1 _04202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14586_ _07754_ _07756_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__xnor2_1
X_11798_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _04910_ vssd1 vssd1 vccd1 vccd1 _04988_
+ sky130_fd_sc_hd__mux2_1
X_19113_ _03142_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__clkbuf_2
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ _08466_ _09184_ _08910_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__a21o_1
XFILLER_119_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13537_ _06682_ _06693_ _06700_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a31o_4
X_10749_ _04143_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__clkbuf_4
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20372__230 clknet_1_0__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__inv_2
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19044_ rbzero.spi_registers.new_other\[4\] _03098_ _03114_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00765_ sky130_fd_sc_hd__o211a_1
X_16256_ _09347_ _09348_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13468_ _06623_ _06627_ _06634_ _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__o211a_2
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15207_ _08290_ _08301_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__or2b_1
X_12419_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _05314_ vssd1 vssd1 vccd1 vccd1 _05604_
+ sky130_fd_sc_hd__mux2_1
X_16187_ _09278_ _09279_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _06540_ _06542_ _06545_ _06553_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__or4_2
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ rbzero.wall_tracer.stepDistY\[-5\] _08157_ _08232_ vssd1 vssd1 vccd1 vccd1
+ _08233_ sky130_fd_sc_hd__o21ai_4
XFILLER_126_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15069_ _08159_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__nor2_2
X_19946_ rbzero.debug_overlay.playerX\[3\] _03559_ _03602_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01179_ sky130_fd_sc_hd__a211o_1
XFILLER_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19877_ net53 rbzero.pov.ss_buffer\[0\] _09734_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__mux2_1
XFILLER_110_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18828_ rbzero.pov.spi_buffer\[23\] rbzero.pov.ready_buffer\[23\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18759_ rbzero.spi_registers.spi_counter\[0\] _02929_ rbzero.spi_registers.spi_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21770_ net296 _01359_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20721_ _08117_ clknet_1_0__leaf__05700_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__and2_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20455__305 clknet_1_0__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__inv_2
X_20652_ _03734_ _03873_ _03875_ _03740_ rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1
+ _01612_ sky130_fd_sc_hd__a32o_1
XFILLER_196_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20583_ _03815_ _03816_ _03812_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a21bo_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21204_ clknet_leaf_10_i_clk _00793_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21135_ clknet_leaf_32_i_clk _00724_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21066_ clknet_leaf_84_i_clk _00655_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20017_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ net50 _05946_ net34 vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__and3_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21968_ net494 _01557_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _04910_ vssd1 vssd1 vccd1 vccd1 _04911_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ clknet_leaf_50_i_clk _00508_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ net425 _01488_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14440_ _06959_ _07423_ _07366_ _07309_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__or4b_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] _04840_ vssd1 vssd1
+ vccd1 vccd1 _04842_ sky130_fd_sc_hd__nor3_1
XFILLER_30_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ _04089_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _06993_ _07360_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__or2_1
X_11583_ _04768_ _04769_ rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a21o_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _09056_ _09058_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__nand2_1
XFILLER_210_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13322_ _06448_ _06467_ _06492_ _06482_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__and4_1
X_17090_ _10109_ _10110_ vssd1 vssd1 vccd1 vccd1 _10111_ sky130_fd_sc_hd__nor2_1
XFILLER_182_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10534_ _03973_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__inv_2
XFILLER_127_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16041_ _09004_ _09128_ _09133_ vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__a21o_1
XFILLER_202_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ rbzero.tex_r1\[32\] rbzero.tex_r1\[33\] _04013_ vssd1 vssd1 vccd1 vccd1 _04015_
+ sky130_fd_sc_hd__mux2_1
X_13253_ _06329_ _06419_ _06421_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__nor4b_1
XFILLER_171_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ rbzero.tex_g1\[8\] _04906_ _05181_ _05389_ _05390_ vssd1 vssd1 vccd1 vccd1
+ _05391_ sky130_fd_sc_hd__a311o_1
XFILLER_182_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13184_ rbzero.wall_tracer.visualWallDist\[-3\] _06327_ _04443_ vssd1 vssd1 vccd1
+ vccd1 _06355_ sky130_fd_sc_hd__a21o_1
X_10396_ _03975_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19800_ rbzero.pov.spi_buffer\[38\] rbzero.pov.spi_buffer\[39\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03511_ sky130_fd_sc_hd__mux2_1
X_12135_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _05010_ vssd1 vssd1 vccd1 vccd1 _05323_
+ sky130_fd_sc_hd__mux2_1
X_17992_ _02187_ _02204_ _02202_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16943_ _09167_ _09677_ vssd1 vssd1 vccd1 vccd1 _09965_ sky130_fd_sc_hd__nor2_1
XFILLER_123_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19731_ rbzero.pov.spi_buffer\[5\] rbzero.pov.spi_buffer\[6\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
X_12066_ rbzero.tex_r1\[53\] _05198_ _05236_ _04939_ vssd1 vssd1 vccd1 vccd1 _05255_
+ sky130_fd_sc_hd__a31o_1
XFILLER_42_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ rbzero.tex_b1\[28\] rbzero.tex_b1\[29\] _04303_ vssd1 vssd1 vccd1 vccd1 _04307_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16874_ _09894_ _09895_ vssd1 vssd1 vccd1 vccd1 _09896_ sky130_fd_sc_hd__nor2_1
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15825_ _08874_ _08877_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__xnor2_1
X_18613_ _02817_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__xnor2_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ _03425_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__clkbuf_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20404__259 clknet_1_0__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__inv_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15756_ _08818_ _08819_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__xnor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ rbzero.debug_overlay.vplaneY\[-9\] vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__inv_2
X_12968_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__clkbuf_4
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14707_ _07806_ _07804_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__and2_1
X_18475_ _02569_ _02685_ _08134_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o21a_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11919_ _05086_ _05093_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nor2_4
X_15687_ _08773_ _08778_ _08781_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__a21oi_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12899_ _06034_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nand2_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _09167_ _01718_ _10342_ _10331_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__o31ai_1
XFILLER_178_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14638_ _07799_ _07801_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17357_ _09822_ _10263_ _10264_ _09812_ _10375_ vssd1 vssd1 vccd1 vccd1 _10376_ sky130_fd_sc_hd__o311a_1
XFILLER_202_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ _07717_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _09396_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__nor2_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17288_ _10305_ _10306_ vssd1 vssd1 vccd1 vccd1 _10307_ sky130_fd_sc_hd__nand2_1
XFILLER_173_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19027_ rbzero.map_overlay.i_otherx\[2\] _03101_ vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__or2_1
X_16239_ _09329_ _09331_ vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__xor2_1
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19929_ rbzero.debug_overlay.playerX\[0\] _08315_ _03582_ vssd1 vssd1 vccd1 vccd1
+ _03589_ sky130_fd_sc_hd__a21o_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21822_ net348 _01411_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21753_ net279 _01342_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20704_ _03914_ _03917_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__and3_1
XFILLER_93_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21684_ clknet_leaf_3_i_clk _01273_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20635_ _03859_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__or2_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21118_ clknet_leaf_71_i_clk _00707_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _07065_ _07085_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__nand2_1
X_21049_ clknet_leaf_73_i_clk _00638_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _07015_ _07041_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__and2_1
XFILLER_41_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15610_ _08700_ _08704_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__xor2_1
X_12822_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] _05997_
+ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nand3_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16590_ rbzero.wall_tracer.stepDistX\[8\] _09426_ _06263_ vssd1 vssd1 vccd1 vccd1
+ _09680_ sky130_fd_sc_hd__mux2_2
XFILLER_62_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ _08404_ _08381_ _08460_ _08456_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__or4_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ net71 _05920_ _05921_ _05055_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__a22o_1
XFILLER_199_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11704_ rbzero.floor_leak\[1\] _04817_ _04893_ rbzero.floor_leak\[0\] vssd1 vssd1
+ vccd1 vccd1 _04894_ sky130_fd_sc_hd__o211a_1
X_18260_ rbzero.spi_registers.new_texadd\[2\]\[19\] rbzero.spi_registers.spi_buffer\[19\]
+ _02478_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ _08555_ _08566_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__xnor2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ net25 _05829_ net26 vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a21o_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17211_ _10228_ _10230_ vssd1 vssd1 vccd1 vccd1 _10231_ sky130_fd_sc_hd__nor2_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14423_ _07316_ _07476_ _07593_ _07592_ _07542_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__o32a_1
X_18191_ _02447_ _02450_ _02448_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__o21a_1
X_11635_ gpout0.hpos\[8\] _04824_ _04420_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a21oi_4
XFILLER_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _08666_ _08382_ _08617_ _09079_ vssd1 vssd1 vccd1 vccd1 _10162_ sky130_fd_sc_hd__or4_1
XFILLER_155_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ _07413_ _07466_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__xor2_2
Xclkbuf_1_1__f__03780_ clknet_0__03780_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03780_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11566_ rbzero.texV\[7\] _04755_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__xor2_1
XFILLER_200_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13305_ _06471_ _06472_ _06411_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a21oi_4
X_10517_ rbzero.tex_r1\[7\] rbzero.tex_r1\[8\] _04035_ vssd1 vssd1 vccd1 vccd1 _04042_
+ sky130_fd_sc_hd__mux2_1
X_17073_ _08950_ _10093_ _09977_ _09691_ vssd1 vssd1 vccd1 vccd1 _10094_ sky130_fd_sc_hd__o211ai_1
XFILLER_144_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14285_ _07431_ _07437_ _07429_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__o21a_1
XFILLER_183_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11497_ gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16024_ _09118_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__buf_2
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13236_ rbzero.wall_tracer.visualWallDist\[3\] _04427_ vssd1 vssd1 vccd1 vccd1 _06407_
+ sky130_fd_sc_hd__or2_1
X_10448_ rbzero.tex_r1\[40\] rbzero.tex_r1\[41\] _04002_ vssd1 vssd1 vccd1 vccd1 _04006_
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _04428_ _06037_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__a21o_1
X_20484__331 clknet_1_0__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__inv_2
XFILLER_151_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12118_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _05305_ vssd1 vssd1 vccd1 vccd1 _05306_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13098_ _06270_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__nor2_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17975_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__and2_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16926_ _09529_ _09653_ _09947_ vssd1 vssd1 vccd1 vccd1 _09948_ sky130_fd_sc_hd__a21boi_1
X_12049_ rbzero.tex_r1\[36\] _04982_ _04924_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16857_ _09873_ _09880_ rbzero.wall_tracer.trackDistX\[-2\] _09879_ vssd1 vssd1 vccd1
+ vccd1 _00537_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _08867_ _08902_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__and2_1
X_16788_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09819_ sky130_fd_sc_hd__nand2_1
X_19576_ _03416_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15739_ _08815_ _08829_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__and2_1
X_18527_ _09764_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18458_ _02673_ _02674_ _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a21o_1
XFILLER_179_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17409_ _01698_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nand2_1
X_18389_ _02618_ _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__and2_1
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22021_ clknet_leaf_53_i_clk _01610_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21805_ net331 _01394_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21736_ net262 _01325_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21667_ clknet_leaf_27_i_clk _01256_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11420_ _04607_ _04608_ _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o21ai_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20618_ _03844_ _03845_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__nand3_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21598_ clknet_leaf_70_i_clk _01187_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11351_ rbzero.spi_registers.texadd0\[19\] _04535_ _04542_ vssd1 vssd1 vccd1 vccd1
+ _04543_ sky130_fd_sc_hd__o21a_1
XFILLER_125_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14070_ _07238_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ rbzero.spi_registers.texadd1\[11\] _04461_ vssd1 vssd1 vccd1 vccd1 _04474_
+ sky130_fd_sc_hd__and2_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13021_ rbzero.wall_tracer.trackDistY\[-4\] vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__inv_2
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17760_ _09528_ _01718_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__or2_1
X_14972_ _08095_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16711_ rbzero.traced_texa\[3\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a22o_1
XFILLER_130_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13923_ _06770_ _06877_ _07093_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__and3_1
X_17691_ _01874_ _01875_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__o21ai_1
XFILLER_208_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19430_ _02481_ rbzero.spi_registers.new_other\[1\] _03338_ vssd1 vssd1 vccd1 vccd1
+ _03340_ sky130_fd_sc_hd__mux2_1
X_16642_ _03971_ _09730_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__nor2_1
X_13854_ _06978_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__and2_1
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ net55 _05945_ _05941_ net52 vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a22o_1
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16573_ _09662_ _09046_ _08816_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__a21oi_1
X_19361_ rbzero.spi_registers.new_vshift\[0\] _03297_ _03299_ _03278_ vssd1 vssd1
+ vccd1 vccd1 _00897_ sky130_fd_sc_hd__o211a_1
XFILLER_16_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _06907_ _06910_ _06908_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__a21oi_1
X_10997_ _04296_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15524_ _08616_ _08618_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__or2_1
XFILLER_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18312_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__nand2_1
XFILLER_31_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12736_ net49 _05910_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a21oi_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ rbzero.spi_registers.new_texadd\[3\]\[13\] _03254_ _03259_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__o211a_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _02496_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
X_15455_ _08151_ _08296_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__nor2_1
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12667_ net25 net24 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nor2_2
XFILLER_163_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14406_ _07531_ _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__nor2_1
X_18174_ _02440_ _02441_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o21ai_1
X_11618_ _04798_ _04800_ _04795_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a21o_1
X_15386_ _08413_ _08414_ _08411_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__a21o_1
XFILLER_128_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12598_ _05774_ _05777_ _05770_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__mux2_1
X_17125_ _10141_ _10142_ _10143_ vssd1 vssd1 vccd1 vccd1 _10145_ sky130_fd_sc_hd__and3_1
X_14337_ _06757_ _07417_ _07366_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__or3_1
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11549_ _04672_ rbzero.map_overlay.i_mapdy\[3\] _04738_ _04653_ vssd1 vssd1 vccd1
+ vccd1 _04739_ sky130_fd_sc_hd__o22a_1
XFILLER_171_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _08816_ _09669_ vssd1 vssd1 vccd1 vccd1 _10077_ sky130_fd_sc_hd__nor2_1
XFILLER_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03794_ _03794_ vssd1 vssd1 vccd1 vccd1 clknet_0__03794_ sky130_fd_sc_hd__clkbuf_16
X_14268_ _07419_ _07427_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__xor2_1
XFILLER_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16007_ rbzero.debug_overlay.playerX\[-6\] vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__clkinv_2
X_13219_ rbzero.wall_tracer.visualWallDist\[-6\] _06062_ _04427_ vssd1 vssd1 vccd1
+ vccd1 _06390_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _07344_ _07369_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__nand2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17958_ _02154_ _02121_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__or2b_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16909_ _09666_ _09674_ vssd1 vssd1 vccd1 vccd1 _09931_ sky130_fd_sc_hd__nand2_1
XFILLER_66_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17889_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__nand2_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19628_ _03447_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19559_ rbzero.spi_registers.new_texadd\[0\]\[21\] rbzero.spi_registers.spi_buffer\[21\]
+ _03380_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
XFILLER_207_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21521_ clknet_leaf_84_i_clk _01110_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21452_ net170 _01041_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21383_ clknet_leaf_21_i_clk _00972_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22004_ net150 _01593_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20196_ rbzero.spi_registers.new_texadd\[3\]\[13\] rbzero.spi_registers.spi_buffer\[13\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XFILLER_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03783_ clknet_0__03783_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03783_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10920_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _04248_ vssd1 vssd1 vccd1 vccd1 _04256_
+ sky130_fd_sc_hd__mux2_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10851_ rbzero.tex_g0\[44\] rbzero.tex_g0\[43\] _04215_ vssd1 vssd1 vccd1 vccd1 _04220_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _06730_ _06726_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__xnor2_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _04183_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ net11 vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__inv_2
XFILLER_185_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21719_ net245 _01308_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ rbzero.wall_tracer.stepDistY\[-9\] _08157_ _08334_ _08161_ vssd1 vssd1 vccd1
+ vccd1 _08335_ sky130_fd_sc_hd__o22ai_4
X_12452_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_61_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _04454_ _04504_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__nand2_1
X_15171_ _08235_ _08246_ _08253_ _08265_ vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__or4_1
XFILLER_197_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12383_ _04826_ _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__or2_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14122_ _07289_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__xnor2_1
X_11334_ _04465_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__buf_4
XFILLER_197_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18930_ rbzero.pov.spi_buffer\[72\] rbzero.pov.ready_buffer\[72\] _02967_ vssd1 vssd1
+ vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
X_14053_ _06710_ _07176_ _07174_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_76_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11265_ rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 _04457_
+ sky130_fd_sc_hd__nor2_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__inv_2
XFILLER_133_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18861_ _02967_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__buf_4
X_11196_ _04400_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17812_ _02044_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18792_ rbzero.pov.spi_buffer\[6\] rbzero.pov.ready_buffer\[6\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
XFILLER_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17743_ _01831_ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__xnor2_2
X_14955_ _04442_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__clkbuf_8
XFILLER_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13906_ _06855_ _06860_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__or2b_1
X_17674_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__or2_1
XFILLER_78_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14886_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19413_ _03330_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16625_ _09583_ _09584_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__nor2_1
XFILLER_165_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13837_ _06957_ _06958_ _06962_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o21a_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _08152_ _08535_ _08409_ _08382_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__or4_1
X_19344_ rbzero.spi_registers.got_new_floor _03288_ vssd1 vssd1 vccd1 vccd1 _03289_
+ sky130_fd_sc_hd__nand2_2
X_13768_ _06935_ _06936_ _06937_ _06938_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15507_ _08573_ _08600_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__and2_1
X_12719_ _05893_ _05896_ _05889_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__mux2_1
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16487_ _09541_ _09577_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19275_ rbzero.spi_registers.new_texadd\[3\]\[6\] _03240_ _03249_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00861_ sky130_fd_sc_hd__o211a_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13699_ _06748_ _06733_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or2_1
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15438_ _08298_ _08340_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__or2_1
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18226_ _02486_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_29_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18157_ _10375_ _02428_ _02364_ rbzero.wall_tracer.trackDistY\[3\] vssd1 vssd1 vccd1
+ vccd1 _00564_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _08011_ _08450_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__or2_1
XFILLER_15_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17108_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _10129_ sky130_fd_sc_hd__or2_1
XFILLER_102_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18088_ _02366_ _02367_ _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17039_ _08166_ _10059_ vssd1 vssd1 vccd1 vccd1 _10060_ sky130_fd_sc_hd__nor2_1
XFILLER_132_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03777_ _03777_ vssd1 vssd1 vccd1 vccd1 clknet_0__03777_ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20050_ _03654_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__clkbuf_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20952_ clknet_leaf_60_i_clk _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ clknet_leaf_44_i_clk _00472_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21504_ clknet_leaf_98_i_clk _01093_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21435_ net153 _01024_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21366_ clknet_leaf_10_i_clk _00955_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21297_ clknet_leaf_30_i_clk _00886_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11050_ rbzero.tex_b1\[12\] rbzero.tex_b1\[13\] _04314_ vssd1 vssd1 vccd1 vccd1 _04324_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20179_ rbzero.spi_registers.new_texadd\[3\]\[5\] rbzero.spi_registers.spi_buffer\[5\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__mux2_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _07908_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__clkbuf_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ rbzero.debug_overlay.facingY\[-8\] _05117_ _05138_ _05140_ vssd1 vssd1 vccd1
+ vccd1 _05141_ sky130_fd_sc_hd__a211o_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_106 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_106/HI zeros[13]
+ sky130_fd_sc_hd__conb_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_117 vssd1 vssd1 vccd1 vccd1 ones[8] top_ew_algofoogle_117/LO sky130_fd_sc_hd__conb_1
X_10903_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _04237_ vssd1 vssd1 vccd1 vccd1 _04247_
+ sky130_fd_sc_hd__mux2_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14671_ _07404_ _07406_ _07832_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__or3b_2
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _05070_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__nand2_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _09371_ _09499_ _09500_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13622_ _06617_ _06792_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__or2_1
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ _04210_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__clkbuf_1
X_17390_ _01673_ _01682_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__xnor2_1
X_16341_ _09432_ _09310_ _06263_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__o21ai_4
XFILLER_38_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _06721_ _06708_ _06723_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__a21o_1
X_10765_ _04174_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19060_ rbzero.map_overlay.i_mapdx\[3\] _03122_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__or2_1
X_12504_ _05662_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__nor2_1
X_16272_ _08304_ _09363_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _06632_ _06631_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__nor2_8
XFILLER_173_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ rbzero.tex_g1\[52\] rbzero.tex_g1\[53\] _04132_ vssd1 vssd1 vccd1 vccd1 _04138_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18011_ _02193_ _02200_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__and2b_1
X_15223_ _08317_ _04692_ _08218_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__mux2_1
X_12435_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _04913_ vssd1 vssd1 vccd1 vccd1 _05620_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15154_ _08143_ _08248_ _08160_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12366_ reg_rgb\[22\] _05551_ _05058_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__mux2_4
XFILLER_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _07259_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__xnor2_1
X_11317_ _04477_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__nand2_1
X_15085_ _06389_ _06362_ _06382_ _08179_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__and4b_1
X_19962_ _08190_ _03611_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__nand2_1
XFILLER_180_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _05481_ _05482_ _04946_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__mux2_1
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14036_ _07154_ _07160_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__or2_1
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18913_ _03038_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03462_ clknet_0__03462_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03462_
+ sky130_fd_sc_hd__clkbuf_16
X_11248_ _04428_ _04435_ _04441_ _04439_ _04442_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a32o_1
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19893_ _03560_ rbzero.pov.ready_buffer\[59\] _03561_ vssd1 vssd1 vccd1 vccd1 _03562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ _03002_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11179_ _04391_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18775_ _02951_ _02963_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__and3_1
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15987_ _09075_ _09081_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ _02014_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__and2b_1
X_14938_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.trackDistX\[2\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08073_ sky130_fd_sc_hd__mux2_1
XFILLER_209_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17657_ _01946_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nor2_1
X_14869_ _06470_ _06575_ _08003_ _07989_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__a31o_1
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _09569_ _09570_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__and2b_1
XFILLER_91_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _01801_ _01876_ _01877_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__and3_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19327_ rbzero.floor_leak\[5\] _03272_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__or2_1
X_16539_ _08731_ _08541_ _09628_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__or3_1
XFILLER_176_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19258_ rbzero.spi_registers.got_new_texadd\[3\] _03096_ vssd1 vssd1 vccd1 vccd1
+ _03239_ sky130_fd_sc_hd__nand2_2
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18209_ rbzero.spi_registers.spi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__buf_4
X_19189_ rbzero.spi_registers.new_texadd\[1\]\[18\] _03188_ _03199_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__o211a_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21220_ clknet_leaf_27_i_clk _00809_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21151_ clknet_leaf_3_i_clk _00740_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20102_ rbzero.pov.ready_buffer\[2\] _03663_ _03705_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01232_ sky130_fd_sc_hd__o211a_1
X_21082_ clknet_leaf_88_i_clk _00671_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20033_ rbzero.pov.ready_buffer\[38\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__and3_1
XFILLER_59_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20267__136 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__inv_2
XFILLER_85_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21984_ net510 _01573_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20935_ clknet_leaf_49_i_clk _00524_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20866_ clknet_leaf_64_i_clk _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20797_ clknet_leaf_47_i_clk _00386_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10550_ _04061_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10481_ rbzero.tex_r1\[24\] rbzero.tex_r1\[25\] _04013_ vssd1 vssd1 vccd1 vccd1 _04023_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12220_ rbzero.tex_g1\[19\] _04910_ _05406_ _04912_ vssd1 vssd1 vccd1 vccd1 _05407_
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21418_ clknet_leaf_2_i_clk _01007_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _05337_ _05338_ _04935_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__mux2_1
XFILLER_151_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21349_ clknet_leaf_35_i_clk _00938_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11102_ _04214_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _04672_ _04704_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or3b_1
X_15910_ _08274_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__clkbuf_4
X_11033_ _04315_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16890_ _09522_ _09649_ _09646_ vssd1 vssd1 vccd1 vccd1 _09912_ sky130_fd_sc_hd__o21ai_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _08919_ _08931_ _08935_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__o21a_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _02769_ _02760_ _02759_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a21oi_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _08812_ _08863_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__xor2_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12984_ _06151_ _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__nor2_2
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17511_ _01801_ _01802_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__nand2_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ rbzero.wall_tracer.stepDistY\[-10\] _07892_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07893_ sky130_fd_sc_hd__mux2_1
X_11935_ rbzero.debug_overlay.vplaneX\[0\] _05115_ _05119_ _05123_ vssd1 vssd1 vccd1
+ vccd1 _05124_ sky130_fd_sc_hd__a211o_1
XFILLER_166_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18491_ _06084_ _06096_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__nand2_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _10345_ _10346_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__nor2_1
XFILLER_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14654_ _06575_ _07813_ _07824_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__o21a_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11866_ _05053_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__nor2_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ _06772_ _06768_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__nor2_1
X_10817_ _04201_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__clkbuf_1
X_17373_ _09525_ _09491_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__or3_1
X_14585_ _07423_ _07444_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__nor2_1
XFILLER_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11797_ _04983_ _04986_ _04937_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__mux2_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19112_ _03140_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__clkbuf_4
X_16324_ _09044_ _09046_ _08434_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__a21oi_1
X_13536_ _06701_ _06702_ _06703_ _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__o211ai_4
X_10748_ _04165_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19043_ rbzero.map_overlay.i_othery\[4\] _03101_ vssd1 vssd1 vccd1 vccd1 _03114_
+ sky130_fd_sc_hd__or2_1
X_16255_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerX\[-4\] _08138_
+ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__mux2_1
X_13467_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__inv_2
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ rbzero.tex_g1\[60\] rbzero.tex_g1\[61\] _04046_ vssd1 vssd1 vccd1 vccd1 _04129_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _08291_ _08299_ _08300_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__a21bo_1
X_12418_ _05601_ _05602_ _05190_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__mux2_1
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16186_ _08370_ _08340_ vssd1 vssd1 vccd1 vccd1 _09279_ sky130_fd_sc_hd__or2_1
XFILLER_86_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13398_ _06485_ _06491_ _06493_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor3_1
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15137_ _07954_ _08147_ _08231_ _08160_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__a211o_1
X_12349_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _04907_ vssd1 vssd1 vccd1 vccd1 _05535_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15068_ rbzero.wall_tracer.stepDistY\[-10\] _08161_ _08162_ vssd1 vssd1 vccd1 vccd1
+ _08163_ sky130_fd_sc_hd__a21o_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19945_ rbzero.pov.ready_buffer\[71\] _03586_ _03600_ _03601_ _03565_ vssd1 vssd1
+ vccd1 vccd1 _03602_ sky130_fd_sc_hd__o221a_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14019_ _07184_ _07189_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19876_ _03550_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18827_ _02993_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18758_ _02952_ _02953_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__nor2_1
XFILLER_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17709_ _01997_ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18689_ _02821_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__inv_2
XFILLER_93_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20720_ _08405_ _03924_ _03930_ _01633_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__o31a_1
XFILLER_169_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20651_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__inv_2
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20582_ _03812_ _03815_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand3b_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__05879_ clknet_0__05879_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05879_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21203_ clknet_leaf_23_i_clk _00792_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21134_ clknet_leaf_27_i_clk _00723_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21065_ clknet_leaf_83_i_clk _00654_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20016_ _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__buf_2
XFILLER_59_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ net493 _01556_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__buf_6
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ clknet_leaf_50_i_clk _00507_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21898_ net424 _01487_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20321__185 clknet_1_1__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__inv_2
XFILLER_70_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ rbzero.row_render.size\[7\] _04840_ rbzero.row_render.size\[8\] vssd1 vssd1
+ vccd1 vccd1 _04841_ sky130_fd_sc_hd__o21a_1
XFILLER_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20849_ clknet_leaf_53_i_clk _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03465_ clknet_0__03465_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03465_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ rbzero.tex_r0\[34\] rbzero.tex_r0\[33\] _04088_ vssd1 vssd1 vccd1 vccd1 _04089_
+ sky130_fd_sc_hd__mux2_1
X_14370_ _07539_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__or2_1
XFILLER_168_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ _04768_ _04770_ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ _06478_ _06479_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__xor2_1
XFILLER_70_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10533_ _04050_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _09004_ _09128_ _09133_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__nand3_1
X_13252_ _06324_ _06328_ _06422_ _06322_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__a31oi_4
XFILLER_196_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10464_ _04014_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12203_ rbzero.tex_g1\[9\] _04905_ _05186_ _04919_ vssd1 vssd1 vccd1 vccd1 _05390_
+ sky130_fd_sc_hd__a31o_1
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _04427_ _06048_ _06052_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__and3_1
XFILLER_159_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10395_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__inv_2
X_12134_ _05320_ _05321_ _04947_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__mux2_1
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17991_ _02188_ _02207_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__xor2_1
XFILLER_124_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19730_ _03474_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
X_16942_ _09955_ _09963_ vssd1 vssd1 vccd1 vccd1 _09964_ sky130_fd_sc_hd__xnor2_2
X_12065_ rbzero.tex_r1\[55\] _04924_ _05253_ _04944_ vssd1 vssd1 vccd1 vccd1 _05254_
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ _04306_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16873_ _09639_ _09892_ _09893_ vssd1 vssd1 vccd1 vccd1 _09895_ sky130_fd_sc_hd__and3_1
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18612_ _02802_ _02804_ _02803_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a21bo_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _08885_ _08918_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__nand2_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ rbzero.spi_registers.new_texadd\[1\]\[13\] rbzero.spi_registers.spi_buffer\[13\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__mux2_1
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18543_ _02745_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__xnor2_1
X_15755_ _08846_ _08848_ _08849_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__a21bo_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12967_ rbzero.map_overlay.i_mapdx\[2\] _06120_ rbzero.map_rom.i_col\[4\] _04720_
+ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a22o_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _05075_ _05080_ _05093_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__nor3_4
X_14706_ _07806_ _07859_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__nor2_1
X_18474_ _02697_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__xnor2_1
X_15686_ _08779_ _08780_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__nand2_1
X_12898_ _06037_ _06041_ _06070_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or4b_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17425_ _10330_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__buf_2
XFILLER_159_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11849_ rbzero.row_render.side _05033_ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14637_ _07796_ _07798_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20296__162 clknet_1_1__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__inv_2
X_17356_ _10373_ _10374_ vssd1 vssd1 vccd1 vccd1 _10375_ sky130_fd_sc_hd__or2_2
XFILLER_147_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14568_ _07723_ _07737_ _07738_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16307_ _08370_ _09397_ _09277_ _09398_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__o31a_1
XFILLER_159_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13519_ _06651_ _06626_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__nor2_1
X_17287_ _10274_ _10304_ vssd1 vssd1 vccd1 vccd1 _10306_ sky130_fd_sc_hd__or2_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14499_ _07642_ _07668_ _07669_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__a21oi_2
X_19026_ rbzero.spi_registers.new_other\[7\] _03098_ _03104_ _03103_ vssd1 vssd1 vccd1
+ vccd1 _00757_ sky130_fd_sc_hd__o211a_1
X_16238_ _09165_ _09210_ _09330_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16169_ _09078_ _09261_ _09134_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19928_ _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__inv_2
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20461__310 clknet_1_1__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__inv_2
X_19859_ rbzero.pov.spi_buffer\[66\] rbzero.pov.spi_buffer\[67\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03542_ sky130_fd_sc_hd__mux2_1
XFILLER_69_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03459_ _03459_ vssd1 vssd1 vccd1 vccd1 clknet_0__03459_ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21821_ net347 _01410_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21752_ net278 _01341_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_opt_3_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20703_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03918_
+ sky130_fd_sc_hd__xnor2_1
X_21683_ clknet_leaf_3_i_clk _01272_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20634_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03860_
+ sky130_fd_sc_hd__and2_1
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21117_ clknet_leaf_71_i_clk _00706_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21048_ clknet_leaf_73_i_clk _00637_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _07017_ _07037_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2_1
XFILLER_90_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15540_ _08578_ _08579_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__xnor2_2
X_12752_ _05916_ _05919_ _05923_ _05929_ _05911_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a32o_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__buf_6
XFILLER_199_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15471_ _08564_ _08565_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__nor2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05861_ _05841_ _05847_ _05851_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__and4bb_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _10076_ _10105_ _10229_ vssd1 vssd1 vccd1 vccd1 _10230_ sky130_fd_sc_hd__a21oi_1
X_14422_ _07542_ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__xnor2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _03972_ _04418_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__or2_1
X_18190_ _02455_ _02456_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__nand2_1
XFILLER_202_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17141_ _08382_ _08618_ _09079_ _08666_ vssd1 vssd1 vccd1 vccd1 _10161_ sky130_fd_sc_hd__o22ai_1
X_14353_ _07473_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__nor2_1
X_11565_ _04753_ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__nand2_1
XFILLER_200_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13304_ _06359_ _06361_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and2_2
X_10516_ _04041_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__clkbuf_1
X_17072_ _10092_ vssd1 vssd1 vccd1 vccd1 _10093_ sky130_fd_sc_hd__buf_2
X_14284_ _07363_ _07454_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__or2_1
X_11496_ rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__inv_2
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13235_ _06398_ _06400_ _06405_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__a21oi_2
X_16023_ _08218_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__clkbuf_4
X_10447_ _04005_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ rbzero.wall_tracer.visualWallDist\[2\] _06327_ _04443_ vssd1 vssd1 vccd1
+ vccd1 _06337_ sky130_fd_sc_hd__a21o_1
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12117_ _05010_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__buf_4
XFILLER_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17974_ _02260_ _02261_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__or2_1
X_13097_ rbzero.wall_tracer.mapY\[8\] _06078_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__nor2_1
X_16925_ _08373_ _09176_ _09651_ vssd1 vssd1 vccd1 vccd1 _09947_ sky130_fd_sc_hd__or3_1
X_12048_ rbzero.tex_r1\[37\] _05198_ _05236_ _04939_ vssd1 vssd1 vccd1 vccd1 _05237_
+ sky130_fd_sc_hd__a31o_1
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19644_ clknet_1_1__leaf__03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__buf_1
X_16856_ _09872_ _09877_ _09878_ _09879_ vssd1 vssd1 vccd1 vccd1 _09880_ sky130_fd_sc_hd__o31a_1
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15807_ _08868_ _08901_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__and2_1
XFILLER_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19575_ rbzero.spi_registers.new_texadd\[1\]\[5\] _02489_ _03383_ vssd1 vssd1 vccd1
+ vccd1 _03416_ sky130_fd_sc_hd__mux2_1
X_16787_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09818_ sky130_fd_sc_hd__or2_1
XFILLER_19_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13999_ _06718_ _06755_ _06738_ _06723_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__o211a_1
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18526_ rbzero.map_rom.i_col\[4\] _09119_ _09776_ vssd1 vssd1 vccd1 vccd1 _02739_
+ sky130_fd_sc_hd__a21oi_1
X_15738_ _08831_ _08832_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__or2_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _02681_ _02670_ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15669_ _08757_ _08763_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__nor2_1
XFILLER_34_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17408_ rbzero.wall_tracer.visualWallDist\[2\] _08421_ _01699_ _01700_ vssd1 vssd1
+ vccd1 vccd1 _01701_ sky130_fd_sc_hd__a31o_1
XFILLER_53_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18388_ _02602_ _02603_ _02619_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a21o_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17339_ _10308_ _10357_ vssd1 vssd1 vccd1 vccd1 _10358_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19009_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ _03084_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22020_ clknet_leaf_49_i_clk _01609_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21804_ net330 _01393_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21735_ net261 _01324_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21666_ clknet_leaf_27_i_clk _01255_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20617_ _03838_ _03842_ _03839_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21597_ clknet_leaf_70_i_clk _01186_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ rbzero.spi_registers.texadd1\[19\] _04461_ _04470_ _04541_ vssd1 vssd1 vccd1
+ vccd1 _04542_ sky130_fd_sc_hd__a211o_1
XFILLER_193_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20433__286 clknet_1_1__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__inv_2
X_11281_ _04464_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__and2_1
X_20479_ clknet_1_1__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__buf_1
X_13020_ rbzero.wall_tracer.trackDistY\[-4\] _06182_ rbzero.wall_tracer.trackDistY\[-5\]
+ _06183_ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__o221a_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14971_ rbzero.wall_tracer.stepDistX\[-9\] _07907_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08095_ sky130_fd_sc_hd__mux2_1
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16710_ rbzero.traced_texa\[2\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__a22o_1
X_13922_ _07091_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__and2_1
X_17690_ _08123_ _01979_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__or3b_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16641_ _04408_ _09729_ vssd1 vssd1 vccd1 vccd1 _09730_ sky130_fd_sc_hd__or2_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13853_ _06726_ _06785_ _06977_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ net39 _05980_ _05946_ _05948_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__and4b_1
X_19360_ rbzero.spi_registers.vshift\[0\] _03298_ vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__or2_1
XFILLER_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16572_ _09044_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10996_ rbzero.tex_b1\[38\] rbzero.tex_b1\[39\] _04292_ vssd1 vssd1 vccd1 vccd1 _04296_
+ sky130_fd_sc_hd__mux2_1
X_13784_ _06947_ _06953_ _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__nand3_1
XFILLER_16_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18311_ _05106_ rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1 vccd1 _02548_
+ sky130_fd_sc_hd__and2_1
XFILLER_71_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15523_ _08617_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__clkbuf_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _05888_ net28 _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__and3_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ rbzero.spi_registers.texadd3\[13\] _03255_ vssd1 vssd1 vccd1 vccd1 _03259_
+ sky130_fd_sc_hd__or2_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ rbzero.spi_registers.new_texadd\[2\]\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
X_15454_ _08165_ _08335_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nor2_1
X_12666_ _05833_ _05822_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11617_ _04795_ _04798_ _04800_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__and3_1
X_14405_ _07551_ _07574_ _07575_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__a21oi_2
XFILLER_129_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18173_ _02434_ _02436_ _02435_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__o21ba_1
X_15385_ _08436_ _08479_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__xnor2_2
XFILLER_128_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12597_ _05775_ _05776_ _05765_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__mux2_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17124_ _10141_ _10142_ _10143_ vssd1 vssd1 vccd1 vccd1 _10144_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14336_ _06982_ _07366_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__or2_1
X_11548_ rbzero.map_overlay.i_mapdy\[0\] vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__inv_2
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _10057_ _10075_ vssd1 vssd1 vccd1 vccd1 _10076_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__03793_ _03793_ vssd1 vssd1 vccd1 vccd1 clknet_0__03793_ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14267_ _07431_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__xor2_1
X_11479_ _04648_ _04667_ rbzero.debug_overlay.playerX\[0\] _04413_ _04668_ vssd1 vssd1
+ vccd1 vccd1 _04669_ sky130_fd_sc_hd__o221a_1
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _09000_ _09100_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__xor2_4
X_13218_ _06387_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__xnor2_2
X_14198_ _07367_ _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__and2_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _06285_ _06287_ _06317_ _06318_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a41o_1
XFILLER_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _02243_ _02244_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__xnor2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16908_ _09650_ _09657_ _09656_ vssd1 vssd1 vccd1 vccd1 _09930_ sky130_fd_sc_hd__a21o_1
X_17888_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__or2_1
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19627_ _03442_ _03443_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and3b_1
X_16839_ _09854_ _09856_ _09855_ vssd1 vssd1 vccd1 vccd1 _09864_ sky130_fd_sc_hd__a21boi_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19558_ _03407_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20222__95 clknet_1_1__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
XFILLER_0_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18509_ _06144_ _09766_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__nor2_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19489_ _03371_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21520_ clknet_leaf_84_i_clk _01109_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21451_ net169 _01040_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21382_ clknet_leaf_28_i_clk _00971_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22003_ net149 _01592_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20195_ _03764_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03782_ clknet_0__03782_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03782_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10850_ _04219_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10781_ rbzero.tex_g1\[12\] rbzero.tex_g1\[13\] _04177_ vssd1 vssd1 vccd1 vccd1 _04183_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _05701_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
X_21718_ net244 _01307_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _05634_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21649_ clknet_leaf_83_i_clk _01238_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_200_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _04590_ _04591_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _06262_ _08257_ _08264_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__o21ai_4
X_12382_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _04893_ vssd1 vssd1 vccd1 vccd1 _05567_
+ sky130_fd_sc_hd__mux2_1
XFILLER_193_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14121_ _07226_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__nor2_1
XFILLER_153_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ _04458_ _04521_ _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__o21ai_1
XFILLER_180_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19685__64 clknet_1_0__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
XFILLER_141_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _07178_ _07222_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13003_ rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__inv_2
X_18860_ _03010_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11195_ rbzero.tex_b0\[8\] rbzero.tex_b0\[7\] _04395_ vssd1 vssd1 vccd1 vccd1 _04400_
+ sky130_fd_sc_hd__mux2_1
X_17811_ _01697_ _09433_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _02974_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ _09542_ _02031_ _01943_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14954_ rbzero.wall_tracer.visualWallDist\[7\] _08046_ vssd1 vssd1 vccd1 vccd1 _08084_
+ sky130_fd_sc_hd__or2_1
XFILLER_169_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _06837_ _07066_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nand2_1
X_17673_ _01771_ _01855_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ _06103_ _08033_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__or2_1
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19412_ _02473_ rbzero.spi_registers.new_leak\[0\] _03329_ vssd1 vssd1 vccd1 vccd1
+ _03330_ sky130_fd_sc_hd__mux2_1
XFILLER_63_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624_ _09610_ _09713_ vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__xnor2_1
X_13836_ _06996_ _07006_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__or2_1
XFILLER_51_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _03096_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__buf_4
X_16555_ _09544_ _09553_ _09644_ vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__a21bo_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10979_ rbzero.tex_b1\[46\] rbzero.tex_b1\[47\] _04281_ vssd1 vssd1 vccd1 vccd1 _04287_
+ sky130_fd_sc_hd__mux2_1
X_13767_ _06935_ _06936_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15506_ _08573_ _08600_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__nor2_1
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12718_ _05894_ _05895_ _05884_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__mux2_1
X_19274_ rbzero.spi_registers.texadd3\[6\] _03242_ vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__or2_1
X_16486_ _09575_ _09576_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__xor2_1
X_13698_ _06700_ _06738_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__nand2_1
X_18225_ rbzero.spi_registers.new_texadd\[2\]\[3\] _02485_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02486_ sky130_fd_sc_hd__mux2_1
X_15437_ _08529_ _08530_ _08329_ _08531_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__a31o_1
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12649_ _05823_ _05825_ _05826_ _05827_ net26 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__a32o_1
XFILLER_89_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18156_ _02341_ _02426_ _02427_ _02339_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__o31a_1
XFILLER_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _08012_ _08450_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__nand2_1
XFILLER_129_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20416__270 clknet_1_1__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__inv_2
XFILLER_172_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17107_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _10128_ sky130_fd_sc_hd__nand2_1
X_14319_ _07316_ _07360_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__or2_1
XFILLER_176_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18087_ _02359_ _02362_ _02360_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__o21ai_1
XFILLER_171_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15299_ _07992_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__xor2_1
XFILLER_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17038_ _08580_ vssd1 vssd1 vccd1 vccd1 _10059_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__03776_ _03776_ vssd1 vssd1 vccd1 vccd1 clknet_0__03776_ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _03079_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__clkbuf_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20951_ clknet_leaf_60_i_clk _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ clknet_leaf_49_i_clk _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21503_ clknet_leaf_82_i_clk _01092_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21434_ net152 _01023_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21365_ clknet_leaf_9_i_clk _00954_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21296_ clknet_leaf_31_i_clk _00885_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20178_ _03755_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20244__115 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__inv_2
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ rbzero.debug_overlay.facingY\[-2\] _05107_ _05122_ rbzero.debug_overlay.facingY\[-9\]
+ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a221o_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_107 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_107/HI zeros[14]
+ sky130_fd_sc_hd__conb_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _04246_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_118 vssd1 vssd1 vccd1 vccd1 ones[9] top_ew_algofoogle_118/LO sky130_fd_sc_hd__conb_1
XFILLER_205_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14670_ _07838_ _07530_ _07802_ _07840_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__o31a_2
X_11882_ _05067_ _05068_ gpout0.hpos\[6\] gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1
+ _05071_ sky130_fd_sc_hd__a2bb2o_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10833_ rbzero.tex_g0\[52\] rbzero.tex_g0\[51\] _04203_ vssd1 vssd1 vccd1 vccd1 _04210_
+ sky130_fd_sc_hd__mux2_1
X_13621_ _06658_ _06783_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16340_ rbzero.trace_state\[0\] rbzero.wall_tracer.stepDistY\[7\] _08338_ vssd1 vssd1
+ vccd1 vccd1 _09432_ sky130_fd_sc_hd__and3_1
X_10764_ rbzero.tex_g1\[20\] rbzero.tex_g1\[21\] _04166_ vssd1 vssd1 vccd1 vccd1 _04174_
+ sky130_fd_sc_hd__mux2_1
X_13552_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__inv_2
XFILLER_197_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ net53 _05659_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a21oi_1
XFILLER_185_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16271_ _09362_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__buf_4
X_13483_ _06651_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__or2_2
XFILLER_200_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10695_ _04137_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18010_ _02212_ _02242_ _02210_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a21o_1
X_12434_ _05617_ _05618_ _04826_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__mux2_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15222_ _08315_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__nand2_1
XFILLER_173_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15153_ _06062_ _06389_ _04463_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__mux2_1
X_12365_ _04661_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__and3b_4
XFILLER_165_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14104_ _07273_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__and2_1
X_11316_ rbzero.texu_hot\[5\] _04476_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__or2_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15084_ rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\] _06375_
+ _06366_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__nor4_1
X_19961_ _08189_ rbzero.pov.ready_buffer\[45\] _03561_ vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12296_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _04908_ vssd1 vssd1 vccd1 vccd1 _05482_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18912_ rbzero.pov.spi_buffer\[63\] rbzero.pov.ready_buffer\[63\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
X_14035_ _06769_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__buf_2
XFILLER_107_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11247_ _04434_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_1_1__f__03461_ clknet_0__03461_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03461_
+ sky130_fd_sc_hd__clkbuf_16
X_19892_ _03437_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__buf_4
XFILLER_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18843_ rbzero.pov.spi_buffer\[30\] rbzero.pov.ready_buffer\[30\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11178_ rbzero.tex_b0\[16\] rbzero.tex_b0\[15\] _04384_ vssd1 vssd1 vccd1 vccd1 _04391_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18774_ rbzero.spi_registers.spi_counter\[6\] _02961_ vssd1 vssd1 vccd1 vccd1 _02964_
+ sky130_fd_sc_hd__nand2_1
XFILLER_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15986_ _09078_ _09080_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__or2_1
X_17725_ _01809_ _01923_ _01925_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a21bo_1
X_14937_ _08065_ _08071_ _08072_ _08061_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__o211a_1
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _01831_ _01945_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__nor2_1
XFILLER_91_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868_ _06568_ _08020_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__or2_1
X_16607_ _09684_ _09696_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__xnor2_1
X_13819_ _06944_ _06940_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__nor2_1
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17587_ _01801_ _01876_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a21oi_2
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14799_ _06581_ _07962_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__or2_1
XFILLER_44_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19326_ rbzero.spi_registers.new_leak\[4\] _03271_ _03277_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00883_ sky130_fd_sc_hd__o211a_1
X_16538_ _08734_ _08617_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__or2_1
XFILLER_17_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19257_ rbzero.spi_registers.new_texadd\[2\]\[23\] _03205_ _03238_ _03237_ vssd1
+ vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__o211a_1
X_16469_ _09559_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__clkbuf_4
XFILLER_149_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18208_ _02329_ _02472_ _02364_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1
+ vccd1 _00571_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_191_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19188_ rbzero.spi_registers.texadd1\[18\] _03189_ vssd1 vssd1 vccd1 vccd1 _03199_
+ sky130_fd_sc_hd__or2_1
XFILLER_145_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19649__31 clknet_1_0__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18139_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] _02409_
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a21o_1
XFILLER_89_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21150_ clknet_leaf_100_i_clk _00739_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19664__45 clknet_1_1__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
X_20101_ rbzero.debug_overlay.vplaneY\[-7\] _03685_ vssd1 vssd1 vccd1 vccd1 _03705_
+ sky130_fd_sc_hd__or2_1
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21081_ clknet_leaf_84_i_clk _00670_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20032_ rbzero.debug_overlay.facingX\[-5\] _03663_ _03666_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01201_ sky130_fd_sc_hd__a211o_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21983_ net509 _01572_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ clknet_leaf_45_i_clk _00523_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ clknet_leaf_65_i_clk _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20796_ clknet_leaf_68_i_clk _00001_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_139_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _04022_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21417_ clknet_leaf_2_i_clk _01006_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12150_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _04948_ vssd1 vssd1 vccd1 vccd1 _05338_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21348_ clknet_leaf_35_i_clk _00937_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _04350_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ _04731_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__and2_1
X_21279_ clknet_leaf_1_i_clk _00868_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ rbzero.tex_b1\[21\] rbzero.tex_b1\[22\] _04314_ vssd1 vssd1 vccd1 vccd1 _04315_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _08932_ _08934_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__nand2_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _08864_ _08865_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__and2_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12983_ _06142_ _06153_ _06156_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__and4bb_2
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _01773_ _01774_ _01800_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__nand3_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14722_ _06633_ _07875_ _07890_ _07891_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__a31o_2
XFILLER_166_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _05120_ _05121_ _05122_ rbzero.debug_overlay.vplaneX\[-9\] vssd1 vssd1 vccd1
+ vccd1 _05123_ sky130_fd_sc_hd__a22o_1
X_18490_ _06086_ _06265_ _02711_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _01726_ _01733_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__xnor2_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14653_ _06574_ _07823_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__nand2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11865_ gpout0.vpos\[8\] _05054_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _05055_
+ sky130_fd_sc_hd__a21o_4
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _06719_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__clkinv_2
X_17372_ _10275_ _01664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__xnor2_1
X_10816_ rbzero.tex_g0\[60\] rbzero.tex_g0\[59\] _04121_ vssd1 vssd1 vccd1 vccd1 _04201_
+ sky130_fd_sc_hd__mux2_1
X_11796_ _04984_ _04985_ _04922_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__mux2_1
XFILLER_186_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14584_ _07417_ _07476_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__nor2_1
X_19111_ rbzero.spi_registers.new_texadd\[0\]\[9\] _03141_ _03154_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00792_ sky130_fd_sc_hd__o211a_1
X_16323_ _09408_ _09414_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ _06655_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__nand2_1
XFILLER_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ rbzero.tex_g1\[28\] rbzero.tex_g1\[29\] _04155_ vssd1 vssd1 vccd1 vccd1 _04165_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19042_ rbzero.spi_registers.new_other\[3\] _03098_ _03113_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00764_ sky130_fd_sc_hd__o211a_1
X_16254_ _09344_ _09346_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__xor2_4
X_10678_ _04128_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__clkbuf_1
X_13466_ _06635_ _06636_ _06589_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__mux2_1
X_15205_ _08245_ _08252_ _08265_ _08275_ vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__or4_1
X_12417_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _05314_ vssd1 vssd1 vccd1 vccd1 _05602_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16185_ _09152_ _09276_ _09277_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__a21o_1
X_13397_ _06537_ _06539_ _06566_ _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__a31o_4
XFILLER_86_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15136_ rbzero.side_hot _06058_ _08142_ _08230_ vssd1 vssd1 vccd1 vccd1 _08231_ sky130_fd_sc_hd__o211a_1
X_12348_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _04907_ vssd1 vssd1 vccd1 vccd1 _05534_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19944_ rbzero.debug_overlay.playerX\[3\] _03594_ _03116_ vssd1 vssd1 vccd1 vccd1
+ _03601_ sky130_fd_sc_hd__a21o_1
X_12279_ _05277_ _05291_ _05465_ _04703_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a31oi_1
X_15067_ rbzero.trace_state\[0\] _06260_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__nor2_8
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _07187_ _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__nor2_1
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19875_ rbzero.pov.mosi rbzero.pov.mosi_buffer\[0\] _03084_ vssd1 vssd1 vccd1 vccd1
+ _03550_ sky130_fd_sc_hd__mux2_1
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20528__371 clknet_1_0__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__inv_2
XFILLER_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18826_ rbzero.pov.spi_buffer\[22\] rbzero.pov.ready_buffer\[22\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02993_ sky130_fd_sc_hd__mux2_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18757_ rbzero.spi_registers.spi_counter\[0\] _02929_ vssd1 vssd1 vccd1 vccd1 _02953_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15969_ _09035_ _09063_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__xnor2_2
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17708_ _10315_ _09243_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__nor2_1
X_18688_ _02821_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02888_
+ sky130_fd_sc_hd__nor2_1
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _01818_ _09677_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__nor2_1
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20650_ _03870_ _03871_ _03872_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__and3_1
XFILLER_143_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ rbzero.spi_registers.new_texadd\[3\]\[21\] _03239_ _03268_ _03265_ vssd1
+ vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__o211a_1
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20581_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03816_
+ sky130_fd_sc_hd__nand2_1
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20273__141 clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__inv_2
XFILLER_178_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21202_ clknet_leaf_22_i_clk _00791_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21133_ clknet_leaf_32_i_clk _00722_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21064_ clknet_leaf_82_i_clk _00653_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20015_ _03095_ _03557_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nand2_1
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ net492 _01555_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ clknet_leaf_50_i_clk _00506_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21897_ net423 _01486_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ rbzero.row_render.size\[6\] _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__and2_1
X_20848_ clknet_leaf_55_i_clk _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03464_ clknet_0__03464_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03464_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20356__216 clknet_1_1__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__inv_2
XFILLER_168_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _04054_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__clkbuf_4
XFILLER_11_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11581_ rbzero.texV\[5\] _04765_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20779_ _03959_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ rbzero.tex_r1\[0\] rbzero.tex_r1\[1\] _04046_ vssd1 vssd1 vccd1 vccd1 _04050_
+ sky130_fd_sc_hd__mux2_1
X_13320_ _06486_ _06487_ _06480_ _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__and4_1
XFILLER_168_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ rbzero.tex_r1\[33\] rbzero.tex_r1\[34\] _04013_ vssd1 vssd1 vccd1 vccd1 _04014_
+ sky130_fd_sc_hd__mux2_1
X_13251_ rbzero.wall_tracer.visualWallDist\[6\] _04427_ vssd1 vssd1 vccd1 vccd1 _06422_
+ sky130_fd_sc_hd__or2_1
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12202_ rbzero.tex_g1\[11\] _04910_ _05388_ _04912_ vssd1 vssd1 vccd1 vccd1 _05389_
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ _06288_ _06347_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__xnor2_2
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__clkbuf_4
XFILLER_151_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12133_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _05010_ vssd1 vssd1 vccd1 vccd1 _05321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _02274_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _09961_ _09962_ vssd1 vssd1 vccd1 vccd1 _09963_ sky130_fd_sc_hd__nand2_1
X_12064_ rbzero.tex_r1\[54\] _05031_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
XFILLER_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11015_ rbzero.tex_b1\[29\] rbzero.tex_b1\[30\] _04303_ vssd1 vssd1 vccd1 vccd1 _04306_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16872_ _09639_ _09892_ _09893_ vssd1 vssd1 vccd1 vccd1 _09894_ sky130_fd_sc_hd__a21oi_4
XFILLER_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18611_ _02800_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__xnor2_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _08879_ _08884_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__or2_1
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19591_ _03424_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__clkbuf_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _05129_ rbzero.wall_tracer.rayAddendY\[-6\] _02753_ vssd1 vssd1 vccd1 vccd1
+ _02754_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _08731_ _08847_ _08473_ _08457_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__or4_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ rbzero.wall_tracer.visualWallDist\[10\] _06137_ _06141_ vssd1 vssd1 vccd1
+ vccd1 _06142_ sky130_fd_sc_hd__or3b_4
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _06575_ _07874_ _06631_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__a21o_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__clkbuf_4
X_18473_ _02598_ rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 _02698_
+ sky130_fd_sc_hd__xnor2_1
X_15685_ _08356_ _08697_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__or2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nand2_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17424_ _10333_ _10334_ _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a21bo_1
XFILLER_166_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _07804_ _07805_ _07806_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__mux2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ rbzero.row_render.side _05037_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__nor2_1
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _10246_ _10254_ _10372_ _08123_ vssd1 vssd1 vccd1 vccd1 _10374_ sky130_fd_sc_hd__a31o_1
XFILLER_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14567_ _07725_ _07736_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nor2_1
X_11779_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _04914_ vssd1 vssd1 vccd1 vccd1 _04969_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _09152_ _09276_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__nand2_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13518_ _06619_ _06622_ _06688_ _06602_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__o211a_1
X_17286_ _10274_ _10304_ vssd1 vssd1 vccd1 vccd1 _10305_ sky130_fd_sc_hd__nand2_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ _07643_ _07667_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__nor2_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ rbzero.map_overlay.i_otherx\[1\] _03101_ vssd1 vssd1 vccd1 vccd1 _03104_
+ sky130_fd_sc_hd__or2_1
X_16237_ _09207_ _09209_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__nor2_1
XFILLER_173_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ _06477_ _06588_ _06578_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__mux2_1
XFILLER_127_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16168_ _09135_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__inv_2
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15119_ _08178_ _08195_ _08201_ _08213_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__o22ai_1
XFILLER_142_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16099_ _08461_ _09053_ _09192_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__nor3_1
XFILLER_141_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19927_ rbzero.debug_overlay.playerX\[0\] _08315_ vssd1 vssd1 vccd1 vccd1 _03587_
+ sky130_fd_sc_hd__or2_1
XFILLER_130_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19858_ _03541_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03458_ _03458_ vssd1 vssd1 vccd1 vccd1 clknet_0__03458_ sky130_fd_sc_hd__clkbuf_16
X_18809_ rbzero.pov.spi_buffer\[14\] rbzero.pov.ready_buffer\[14\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02984_ sky130_fd_sc_hd__mux2_1
X_19789_ _03505_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21820_ net346 _01409_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21751_ net277 _01340_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20702_ _09732_ _03916_ _03917_ _03740_ rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1
+ _01620_ sky130_fd_sc_hd__a32o_1
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21682_ clknet_leaf_100_i_clk _01271_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20633_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__nor2_1
XFILLER_20_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21116_ clknet_leaf_13_i_clk _00705_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21047_ clknet_leaf_87_i_clk _00636_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand2_1
XFILLER_189_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__04634_ clknet_0__04634_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04634_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _05884_ _05889_ _05925_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__a31o_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ net475 _01538_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11702_ _04785_ _04828_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__nand2_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15470_ _08561_ _08563_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__and2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05711_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__clkinv_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _07591_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__inv_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11633_ _04806_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nor2_8
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17140_ _10043_ _10046_ _10044_ vssd1 vssd1 vccd1 vccd1 _10160_ sky130_fd_sc_hd__a21bo_1
XFILLER_168_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14352_ _07475_ _07518_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__o21a_1
XFILLER_196_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11564_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _04754_ sky130_fd_sc_hd__or2_1
XFILLER_11_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _06471_ _06473_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__xnor2_4
X_10515_ rbzero.tex_r1\[8\] rbzero.tex_r1\[9\] _04035_ vssd1 vssd1 vccd1 vccd1 _04041_
+ sky130_fd_sc_hd__mux2_1
X_17071_ _09970_ _09972_ vssd1 vssd1 vccd1 vccd1 _10092_ sky130_fd_sc_hd__and2_1
XFILLER_196_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14283_ _07448_ _07449_ _07453_ _07211_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__o2bb2a_1
X_11495_ gpout0.vpos\[1\] rbzero.debug_overlay.playerY\[-2\] vssd1 vssd1 vccd1 vccd1
+ _04685_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ _09104_ _09116_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10446_ rbzero.tex_r1\[41\] rbzero.tex_r1\[42\] _04002_ vssd1 vssd1 vccd1 vccd1 _04005_
+ sky130_fd_sc_hd__mux2_1
X_13234_ _04444_ _06402_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__a21oi_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _04444_ _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__nand2_1
XFILLER_3_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20410__265 clknet_1_1__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__inv_2
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ _04906_ _05301_ _05303_ _04920_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__o211a_1
X_17973_ _02169_ _02173_ _02259_ _01757_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a31o_1
X_13096_ rbzero.wall_tracer.mapY\[8\] _06078_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__and2_1
XFILLER_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16924_ _09944_ _09945_ vssd1 vssd1 vccd1 vccd1 _09946_ sky130_fd_sc_hd__xor2_1
X_12047_ _04829_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19643_ clknet_1_0__leaf__04634_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__buf_1
X_16855_ _09782_ vssd1 vssd1 vccd1 vccd1 _09879_ sky130_fd_sc_hd__buf_4
XFILLER_20_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15806_ _08900_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__inv_2
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19574_ _03415_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__clkbuf_1
X_16786_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ _09810_ vssd1 vssd1 vccd1 vccd1 _09817_ sky130_fd_sc_hd__a21o_1
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13998_ _06721_ _06758_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__nand2_1
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18525_ _02738_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
X_15737_ _08804_ _08801_ _08803_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__a21oi_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ rbzero.wall_tracer.mapY\[6\] rbzero.wall_tracer.mapY\[9\] rbzero.wall_tracer.mapY\[8\]
+ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or4_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _02598_ _02569_ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a21oi_1
X_15668_ _08761_ _08762_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__or2_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20339__200 clknet_1_1__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__inv_2
XFILLER_178_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _01697_ _09044_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__nor2_1
XFILLER_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14619_ _07745_ _07788_ _07789_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__a21o_1
X_18387_ _02592_ _02602_ _02588_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__o21a_1
X_20491__337 clknet_1_0__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__inv_2
X_15599_ _08680_ _08692_ _08693_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17338_ _10355_ _10356_ vssd1 vssd1 vccd1 vccd1 _10357_ sky130_fd_sc_hd__nor2_1
XFILLER_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ rbzero.wall_tracer.visualWallDist\[2\] _08421_ vssd1 vssd1 vccd1 vccd1 _10288_
+ sky130_fd_sc_hd__nand2_2
XFILLER_174_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19008_ _03089_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20385__242 clknet_1_1__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__inv_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21803_ net329 _01392_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ net260 _01323_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21665_ clknet_leaf_27_i_clk _01254_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20616_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__nand2_1
XFILLER_177_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21596_ clknet_leaf_69_i_clk _01185_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ rbzero.spi_registers.texadd0\[12\] _04467_ _04468_ _04471_ vssd1 vssd1 vccd1
+ vccd1 _04472_ sky130_fd_sc_hd__o22a_1
XFILLER_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19700__77 clknet_1_0__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14970_ _08094_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13921_ _07089_ _07090_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__or2_1
XFILLER_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16640_ _09728_ vssd1 vssd1 vccd1 vccd1 _09729_ sky130_fd_sc_hd__clkbuf_4
X_13852_ _07021_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _05976_ _05977_ _05978_ _05979_ net38 vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__a32o_1
X_16571_ _09643_ _09660_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13783_ _06949_ _06950_ _06952_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__a21o_1
X_10995_ _04295_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18310_ _05106_ rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__nor2_1
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15522_ rbzero.wall_tracer.visualWallDist\[4\] _08149_ vssd1 vssd1 vccd1 vccd1 _08617_
+ sky130_fd_sc_hd__nand2_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _05711_ _05911_ net50 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21o_1
XFILLER_31_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19290_ rbzero.spi_registers.new_texadd\[3\]\[12\] _03254_ _03258_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__o211a_1
XFILLER_71_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18241_ _02495_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15453_ _08524_ _08520_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__or2b_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _05055_ _05842_ _05843_ net71 vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a22oi_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14404_ _07552_ _07573_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__nor2_1
X_18172_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__and2_1
X_11616_ _04802_ _04804_ _04805_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__o21a_4
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15384_ _08469_ _08478_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__xor2_2
XFILLER_204_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12596_ _03975_ _04420_ _05763_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__mux2_1
XFILLER_184_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17123_ _10035_ _10037_ _10038_ _10039_ vssd1 vssd1 vccd1 vccd1 _10143_ sky130_fd_sc_hd__o22a_1
XFILLER_117_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14335_ _07423_ _07303_ _07398_ _06959_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__o22a_1
X_11547_ rbzero.map_overlay.i_mapdy\[5\] _04736_ _04670_ vssd1 vssd1 vccd1 vccd1 _04737_
+ sky130_fd_sc_hd__o21a_1
XFILLER_204_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17054_ _10058_ _10074_ vssd1 vssd1 vccd1 vccd1 _10075_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03792_ _03792_ vssd1 vssd1 vccd1 vccd1 clknet_0__03792_ sky130_fd_sc_hd__clkbuf_16
X_14266_ _06993_ _07249_ _07432_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__o31a_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11478_ _04651_ rbzero.debug_overlay.playerY\[1\] vssd1 vssd1 vccd1 vccd1 _04668_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ _09098_ _09099_ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__and2_2
X_20334__196 clknet_1_0__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__inv_2
X_13217_ _06297_ _06304_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__and2b_1
X_10429_ rbzero.tex_r1\[49\] rbzero.tex_r1\[50\] _03991_ vssd1 vssd1 vccd1 vccd1 _03996_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14197_ _07253_ _07045_ _07366_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13148_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__nor2_1
XFILLER_97_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17956_ _02118_ _02119_ _02156_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__o21a_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _06249_ _06252_ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__o21ai_2
X_16907_ _09897_ _09928_ vssd1 vssd1 vccd1 vccd1 _09929_ sky130_fd_sc_hd__xnor2_1
X_17887_ _02173_ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nand2_1
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19626_ _03439_ _03445_ _03440_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__a21boi_1
XFILLER_66_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16838_ _09861_ _09862_ vssd1 vssd1 vccd1 vccd1 _09863_ sky130_fd_sc_hd__or2b_1
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19557_ rbzero.spi_registers.new_texadd\[0\]\[20\] rbzero.spi_registers.spi_buffer\[20\]
+ _03380_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ _09784_ _09801_ _09802_ _09785_ rbzero.wall_tracer.mapX\[10\] vssd1 vssd1
+ vccd1 vccd1 _00527_ sky130_fd_sc_hd__a32o_1
XFILLER_20_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18508_ _02725_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19488_ rbzero.spi_registers.new_mapd\[8\] rbzero.spi_registers.spi_buffer\[8\] _03362_
+ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__mux2_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18439_ _02664_ _02665_ _02662_ _02663_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o211ai_2
XFILLER_210_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21450_ net168 _01039_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ clknet_1_0__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__buf_1
X_21381_ clknet_leaf_28_i_clk _00970_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22002_ net148 _01591_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20194_ rbzero.spi_registers.new_texadd\[3\]\[12\] rbzero.spi_registers.spi_buffer\[12\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__mux2_1
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03781_ clknet_0__03781_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03781_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _04182_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21717_ net243 _01306_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ reg_vsync _04431_ _05058_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__mux2_2
X_21648_ clknet_leaf_83_i_clk _01237_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _04506_ _04485_ _04504_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a31o_1
X_12381_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _04931_ vssd1 vssd1 vccd1 vccd1 _05566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21579_ clknet_leaf_70_i_clk _01168_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_181_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14120_ _07264_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__xnor2_1
X_11332_ rbzero.spi_registers.texadd0\[15\] _04467_ _04523_ vssd1 vssd1 vccd1 vccd1
+ _04524_ sky130_fd_sc_hd__o21a_1
XFILLER_192_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14051_ _07220_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nand2_1
X_11263_ rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 _04455_
+ sky130_fd_sc_hd__and2_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _06174_ _06176_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__or3b_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ _04399_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17810_ _02098_ _02034_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__nand2_1
X_18790_ rbzero.pov.spi_buffer\[5\] rbzero.pov.ready_buffer\[5\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_121_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17741_ _09542_ _10093_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__nor2_1
XFILLER_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14953_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.trackDistX\[7\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__mux2_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13904_ _06868_ _06871_ _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__o21ai_2
X_17672_ _01852_ _01854_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nor2_1
XFILLER_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14884_ _06160_ _06257_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__nand2_4
XFILLER_208_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20522__366 clknet_1_0__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__inv_2
X_16623_ _09711_ _09712_ vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__xor2_1
X_19411_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__buf_2
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13835_ _07002_ _07004_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16554_ _09546_ _09552_ vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__nand2_1
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ rbzero.spi_registers.new_sky\[5\] _03280_ _03287_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00890_ sky130_fd_sc_hd__o211a_1
X_13766_ _06728_ _06807_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nand2_1
X_10978_ _04286_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _08592_ _08598_ _08599_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__a21boi_1
X_12717_ _03975_ _04420_ net28 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__mux2_1
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19273_ rbzero.spi_registers.new_texadd\[3\]\[5\] _03240_ _03248_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00860_ sky130_fd_sc_hd__o211a_1
X_16485_ _09415_ _09443_ _09442_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__a21boi_2
XFILLER_149_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13697_ _06728_ _06758_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__nand2_1
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ rbzero.spi_registers.spi_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__buf_4
X_15436_ _08253_ _08328_ _08325_ _08276_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__o22a_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _05382_ _05470_ _05551_ _05632_ _05822_ net25 vssd1 vssd1 vccd1 vccd1 _05827_
+ sky130_fd_sc_hd__mux4_1
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18155_ _02417_ _02421_ _02424_ _02425_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a211oi_2
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15367_ rbzero.wall_tracer.stepDistY\[4\] _08405_ vssd1 vssd1 vccd1 vccd1 _08462_
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12579_ _05470_ _05719_ _05721_ _05713_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__and4b_1
XFILLER_184_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17106_ _09822_ _10126_ vssd1 vssd1 vccd1 vccd1 _10127_ sky130_fd_sc_hd__nand2_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ _06993_ _07208_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__or2_1
X_18086_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__nand2_1
XFILLER_172_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15298_ _06516_ _07975_ _07981_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__or3b_2
X_17037_ _09955_ _09962_ _09961_ vssd1 vssd1 vccd1 vccd1 _10058_ sky130_fd_sc_hd__a21bo_1
X_14249_ _06854_ _07309_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__and2_1
XFILLER_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ rbzero.spi_registers.spi_cmd\[0\] rbzero.spi_registers.mosi _03078_ vssd1
+ vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _02044_ _02100_ _02102_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a21bo_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20950_ clknet_leaf_59_i_clk _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19609_ _03433_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20881_ clknet_leaf_53_i_clk _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_20497__343 clknet_1_1__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__inv_2
XFILLER_183_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21502_ clknet_leaf_98_i_clk _01091_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21433_ net151 _01022_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21364_ clknet_leaf_22_i_clk _00953_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21295_ clknet_leaf_35_i_clk _00884_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20246_ clknet_1_0__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__buf_1
XFILLER_157_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20177_ rbzero.spi_registers.new_texadd\[3\]\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__mux2_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ rbzero.debug_overlay.facingY\[-5\] _05112_ _05113_ rbzero.debug_overlay.facingY\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a22o_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ rbzero.tex_g0\[20\] rbzero.tex_g0\[19\] _04237_ vssd1 vssd1 vccd1 vccd1 _04246_
+ sky130_fd_sc_hd__mux2_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_108 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_108/HI zeros[15]
+ sky130_fd_sc_hd__conb_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_119 vssd1 vssd1 vccd1 vccd1 ones[10] top_ew_algofoogle_119/LO sky130_fd_sc_hd__conb_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11881_ _05067_ _05068_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or3_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ _06790_ _06717_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__or2_1
XFILLER_38_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10832_ _04209_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ _06617_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__buf_2
X_10763_ _04173_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net52 _05637_ _05664_ net55 vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__a22o_1
X_16270_ rbzero.wall_tracer.visualWallDist\[8\] _08475_ vssd1 vssd1 vccd1 vccd1 _09362_
+ sky130_fd_sc_hd__nand2_4
X_13482_ _06624_ _06652_ _06576_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__mux2_1
XFILLER_185_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10694_ rbzero.tex_g1\[53\] rbzero.tex_g1\[54\] _04132_ vssd1 vssd1 vccd1 vccd1 _04137_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15221_ rbzero.debug_overlay.playerX\[-2\] _08277_ rbzero.debug_overlay.playerX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__o21ai_1
X_12433_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _04893_ vssd1 vssd1 vccd1 vccd1 _05618_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15152_ _07891_ _07942_ _07943_ _08147_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__o31ai_2
X_12364_ _05051_ _05056_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__and2_1
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14103_ _07266_ _07272_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__nand2_1
X_11315_ _04485_ _04504_ _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a21o_1
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ rbzero.wall_tracer.stepDistX\[-3\] _06262_ _08177_ vssd1 vssd1 vccd1 vccd1
+ _08178_ sky130_fd_sc_hd__o21bai_4
X_19960_ _03611_ _03612_ _03613_ _03579_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__o211a_1
X_12295_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _05009_ vssd1 vssd1 vccd1 vccd1 _05481_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18911_ _03037_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
X_14034_ _06720_ _07204_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__03460_ clknet_0__03460_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03460_
+ sky130_fd_sc_hd__clkbuf_16
X_11246_ _04439_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__nor2_1
X_19891_ rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__inv_2
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18842_ _03001_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
X_11177_ _04390_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15985_ _08304_ _08618_ _09079_ _08616_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__o22a_1
X_18773_ rbzero.spi_registers.spi_counter\[6\] _02961_ vssd1 vssd1 vccd1 vccd1 _02963_
+ sky130_fd_sc_hd__or2_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17724_ _02011_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__xor2_1
X_14936_ rbzero.wall_tracer.visualWallDist\[1\] _08046_ vssd1 vssd1 vccd1 vccd1 _08072_
+ sky130_fd_sc_hd__or2_1
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17655_ _01831_ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__and2_1
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ _07826_ _07977_ _07978_ _07979_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__a31o_1
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16606_ _09693_ _09695_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__xor2_1
X_13818_ _06986_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__and2_1
XFILLER_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17586_ _01780_ _01781_ _01782_ _01783_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__o22a_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ _06574_ _07959_ _07960_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__o31a_1
XFILLER_32_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ _09520_ _08541_ _08618_ _09525_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__o22a_1
XFILLER_177_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19325_ _03212_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__clkbuf_4
X_13749_ _06906_ _06916_ _06918_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__or3_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16468_ rbzero.wall_tracer.stepDistX\[7\] _09045_ _09433_ vssd1 vssd1 vccd1 vccd1
+ _09559_ sky130_fd_sc_hd__a21boi_4
X_19256_ rbzero.spi_registers.texadd2\[23\] _03207_ vssd1 vssd1 vccd1 vccd1 _03238_
+ sky130_fd_sc_hd__or2_1
XFILLER_148_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15419_ _08505_ _08513_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__and2_1
X_18207_ _09872_ _02471_ _02337_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__o21a_1
X_19187_ rbzero.spi_registers.new_texadd\[1\]\[17\] _03188_ _03198_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__o211a_1
XFILLER_157_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16399_ rbzero.wall_tracer.visualWallDist\[9\] _08475_ vssd1 vssd1 vccd1 vccd1 _09490_
+ sky130_fd_sc_hd__nand2_2
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18138_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__or2_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18069_ _09823_ _02352_ _02340_ rbzero.wall_tracer.trackDistY\[-9\] vssd1 vssd1 vccd1
+ vccd1 _00552_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20100_ rbzero.pov.ready_buffer\[1\] _03684_ _03704_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01231_ sky130_fd_sc_hd__o211a_1
X_21080_ clknet_leaf_84_i_clk _00669_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20031_ rbzero.pov.ready_buffer\[37\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__and3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20505__350 clknet_1_0__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__inv_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21982_ net508 _01571_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20933_ clknet_leaf_20_i_clk _00522_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_54_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ clknet_leaf_65_i_clk _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20795_ clknet_leaf_68_i_clk _00000_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_168_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21416_ clknet_leaf_1_i_clk _01005_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21347_ clknet_leaf_35_i_clk _00936_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20250__120 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__inv_2
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _04340_ vssd1 vssd1 vccd1 vccd1 _04350_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ gpout0.vpos\[7\] _04653_ _03972_ _04410_ vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__or4_1
XFILLER_150_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21278_ clknet_leaf_1_i_clk _00867_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11031_ _04143_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ _08765_ _08808_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__xor2_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12982_ rbzero.map_rom.b6 rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\] _06157_ vssd1
+ vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__or4_1
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14721_ _06516_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__clkbuf_4
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11933_ _05086_ _05116_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__nor2_4
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _01731_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nor2_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14652_ _07816_ _07821_ _07822_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ gpout0.vpos\[7\] _04648_ _04656_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and3_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13603_ _06770_ _06773_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__nand2_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _09519_ _09242_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nor2_1
X_10815_ _04200_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__clkbuf_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14583_ _06959_ _07361_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__or2_1
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11795_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _04978_ vssd1 vssd1 vccd1 vccd1 _04985_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16322_ _09409_ _09413_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__xnor2_1
X_19110_ rbzero.spi_registers.texadd0\[9\] _03143_ vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__or2_1
XFILLER_186_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13534_ _06680_ _06704_ _06594_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__mux2_1
X_10746_ _04164_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19041_ rbzero.map_overlay.i_othery\[3\] _03101_ vssd1 vssd1 vccd1 vccd1 _03113_
+ sky130_fd_sc_hd__or2_1
X_16253_ _09000_ _09100_ _09226_ _09345_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__a31o_4
XFILLER_51_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13465_ _06506_ _06555_ _06578_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__mux2_1
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ rbzero.tex_g1\[61\] rbzero.tex_g1\[62\] _04046_ vssd1 vssd1 vccd1 vccd1 _04128_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15204_ _08287_ _08298_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12416_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _05314_ vssd1 vssd1 vccd1 vccd1 _05601_
+ sky130_fd_sc_hd__mux2_1
X_16184_ _08368_ _08327_ _08384_ _08813_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__o22a_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13396_ _06486_ _06541_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__nor2_2
XFILLER_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15135_ rbzero.side_hot _06362_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__nand2_1
X_12347_ _05198_ _05532_ _04939_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__o21a_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19943_ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__inv_2
X_15066_ _08160_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__clkbuf_8
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12278_ _04741_ _05292_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__nor2_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _07133_ _07186_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__and2_1
X_11229_ _04051_ _04419_ _04420_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and4_1
X_19874_ _03549_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18825_ _02992_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ _02929_ _02950_ _02951_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a21bo_1
XFILLER_209_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15968_ _09060_ _09062_ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__xnor2_2
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17707_ _08404_ _09363_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__nor2_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14919_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.trackDistX\[-3\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__mux2_1
XFILLER_209_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15899_ _08810_ _08866_ _08991_ _08993_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__a22o_2
X_18687_ _02821_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02887_
+ sky130_fd_sc_hd__and2_1
X_17638_ _01814_ _01928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _10383_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19308_ rbzero.spi_registers.texadd3\[21\] _03241_ vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__or2_1
X_20580_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03815_
+ sky130_fd_sc_hd__or2_1
XFILLER_210_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19239_ rbzero.spi_registers.texadd2\[15\] _03222_ vssd1 vssd1 vccd1 vccd1 _03229_
+ sky130_fd_sc_hd__or2_1
XFILLER_143_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21201_ clknet_leaf_21_i_clk _00790_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21132_ clknet_leaf_29_i_clk _00721_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21063_ clknet_leaf_82_i_clk _00652_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20014_ _03651_ _03653_ _03103_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__o21a_1
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ net491 _01554_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ clknet_leaf_48_i_clk _00505_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21896_ net422 _01485_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20847_ clknet_leaf_57_i_clk _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03463_ clknet_0__03463_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03463_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10600_ _04087_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ rbzero.texV\[4\] _04768_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__nand3_1
X_20778_ _03728_ _03957_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__and3_1
XFILLER_156_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _04049_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _06324_ _06328_ _06420_ _06322_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a31o_1
XFILLER_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ _03979_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12201_ rbzero.tex_g1\[10\] _05236_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or2_1
XFILLER_170_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _04427_ _06071_ _06072_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a31o_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10393_ net47 net48 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__xor2_4
XFILLER_191_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _04964_ vssd1 vssd1 vccd1 vccd1 _05320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16940_ _09956_ _09960_ vssd1 vssd1 vccd1 vccd1 _09962_ sky130_fd_sc_hd__or2_1
X_12063_ rbzero.tex_r1\[56\] _04935_ _04933_ _05250_ _05251_ vssd1 vssd1 vccd1 vccd1
+ _05252_ sky130_fd_sc_hd__a311o_1
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _04305_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16871_ _09620_ _09622_ _09618_ _09619_ vssd1 vssd1 vccd1 vccd1 _09893_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18610_ _02814_ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__nor2_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _08887_ _08892_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__xnor2_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ rbzero.spi_registers.new_texadd\[1\]\[12\] rbzero.spi_registers.spi_buffer\[12\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__mux2_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _08731_ _08473_ _08457_ _08847_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__o22ai_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18541_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] _02752_
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a21o_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12965_ rbzero.wall_tracer.visualWallDist\[9\] rbzero.wall_tracer.visualWallDist\[8\]
+ _06138_ _06140_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__or4_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _05073_ _05091_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a21o_2
X_14704_ _07871_ _07873_ _06580_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__mux2_1
X_15684_ _08356_ _08697_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__nand2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _02688_ _02692_ _02689_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a21bo_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _05999_ _06020_ _06048_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__nand3_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _09542_ _09677_ _10335_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__or3_1
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14635_ _06579_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__buf_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11847_ rbzero.row_render.texu\[0\] _04818_ _05031_ _05036_ vssd1 vssd1 vccd1 vccd1
+ _05037_ sky130_fd_sc_hd__o31ai_2
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _10246_ _10254_ _10372_ vssd1 vssd1 vccd1 vccd1 _10373_ sky130_fd_sc_hd__a21oi_1
X_14566_ _07725_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__xor2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _04920_ _04961_ _04966_ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__a211o_1
X_16305_ _08535_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__clkbuf_4
X_19706__83 clknet_1_1__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13517_ _06643_ _06647_ _06648_ _06598_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a22oi_1
X_17285_ _10286_ _10303_ vssd1 vssd1 vccd1 vccd1 _10304_ sky130_fd_sc_hd__xor2_1
X_10729_ rbzero.tex_g1\[37\] rbzero.tex_g1\[38\] _04155_ vssd1 vssd1 vccd1 vccd1 _04156_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _07643_ _07667_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__xor2_1
X_16236_ _09288_ _09328_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__xnor2_2
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19024_ rbzero.spi_registers.new_other\[6\] _03098_ _03102_ _03103_ vssd1 vssd1 vccd1
+ vccd1 _00756_ sky130_fd_sc_hd__o211a_1
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__buf_2
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16167_ _09247_ _09259_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13379_ _06458_ _06465_ _06531_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or3b_1
XFILLER_138_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15118_ _08212_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__buf_2
XFILLER_142_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ _08042_ _08338_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__or3_2
XFILLER_173_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19926_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__buf_2
X_15049_ _08143_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_74_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19857_ rbzero.pov.spi_buffer\[65\] rbzero.pov.spi_buffer\[66\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03541_ sky130_fd_sc_hd__mux2_1
XFILLER_69_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03457_ _03457_ vssd1 vssd1 vccd1 vccd1 clknet_0__03457_ sky130_fd_sc_hd__clkbuf_16
X_18808_ _02983_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19788_ rbzero.pov.spi_buffer\[32\] rbzero.pov.spi_buffer\[33\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03505_ sky130_fd_sc_hd__mux2_1
XFILLER_209_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_89_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18739_ _02931_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nand2_1
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21750_ net276 _01339_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20701_ _03908_ _03913_ _03914_ _03915_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nand4_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21681_ clknet_leaf_100_i_clk _01270_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20632_ _03734_ _03857_ _03858_ _03740_ rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1
+ _01609_ sky130_fd_sc_hd__a32o_1
XFILLER_20_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21115_ clknet_leaf_13_i_clk _00704_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__05820_ clknet_0__05820_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05820_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21046_ clknet_leaf_87_i_clk _00635_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20362__221 clknet_1_0__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__inv_2
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12750_ clknet_1_0__leaf__04634_ _05910_ _05909_ _05927_ vssd1 vssd1 vccd1 vccd1
+ _05928_ sky130_fd_sc_hd__a31o_2
X_21948_ net474 _01537_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ _04817_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__buf_4
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12681_ _05832_ _05840_ _05859_ net26 vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__o22ai_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ net405 _01468_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14420_ _07306_ _07443_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__nor2_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20561__21 clknet_1_1__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
X_11632_ _04793_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__xnor2_4
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _07519_ _07521_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__or2b_1
X_11563_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _04753_ sky130_fd_sc_hd__nand2_1
XFILLER_7_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _06411_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nor2_2
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10514_ _04040_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__clkbuf_1
X_17070_ _10088_ _10090_ vssd1 vssd1 vccd1 vccd1 _10091_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14282_ _07206_ _07209_ _07205_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__o21a_1
XFILLER_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ rbzero.debug_overlay.playerX\[-3\] _03969_ vssd1 vssd1 vccd1 vccd1 _04684_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_171_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16021_ _09107_ _09114_ _09115_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__a21o_1
X_13233_ _06327_ _06043_ _06054_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__o31a_1
XFILLER_196_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10445_ _04004_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13164_ _06320_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__xnor2_2
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ _05191_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__or2_1
XFILLER_112_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17972_ _02169_ _02173_ _02259_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a21oi_1
X_13095_ rbzero.wall_tracer.mapY\[7\] _06265_ _06266_ _06269_ vssd1 vssd1 vccd1 vccd1
+ _00387_ sky130_fd_sc_hd__a22o_1
XFILLER_123_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19711_ clknet_1_0__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__buf_1
X_16923_ _09397_ _08497_ vssd1 vssd1 vccd1 vccd1 _09945_ sky130_fd_sc_hd__nor2_1
X_12046_ rbzero.tex_r1\[39\] _04924_ _05234_ _04944_ vssd1 vssd1 vccd1 vccd1 _05235_
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19642_ rbzero.pov.spi_counter\[6\] _03454_ _03456_ vssd1 vssd1 vccd1 vccd1 _01021_
+ sky130_fd_sc_hd__o21a_1
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16854_ _09874_ _09875_ _09876_ vssd1 vssd1 vccd1 vccd1 _09878_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _08895_ _08898_ _08899_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__a21o_1
X_19573_ rbzero.spi_registers.new_texadd\[1\]\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__mux2_1
XFILLER_207_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16785_ _06188_ _09786_ _09816_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13997_ _07114_ _07129_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__a21o_1
XFILLER_168_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18524_ rbzero.map_rom.i_col\[4\] _02737_ _09844_ vssd1 vssd1 vccd1 vccd1 _02738_
+ sky130_fd_sc_hd__mux2_1
X_15736_ _08804_ _08801_ _08803_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__and3_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _06110_ _06116_ _06119_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or4_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18455_ _02569_ rbzero.debug_overlay.vplaneX\[-1\] _02598_ vssd1 vssd1 vccd1 vccd1
+ _02682_ sky130_fd_sc_hd__a21oi_1
XFILLER_209_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15667_ _08758_ _08760_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__and2_1
X_12879_ _06043_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nor2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _08475_ _08445_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__and2_1
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _07714_ _07744_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__and2_1
X_15598_ _08663_ _08679_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__nor2_1
X_18386_ _02616_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__and2b_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17337_ _10352_ _10354_ vssd1 vssd1 vccd1 vccd1 _10356_ sky130_fd_sc_hd__and2_1
XFILLER_193_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14549_ _07675_ _07718_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__or2_1
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17268_ _10161_ _10164_ _10162_ vssd1 vssd1 vccd1 vccd1 _10287_ sky130_fd_sc_hd__a21bo_1
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19007_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[0\]
+ _03084_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
XFILLER_162_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16219_ _09192_ _09311_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17199_ _10216_ _10218_ vssd1 vssd1 vccd1 vccd1 _10219_ sky130_fd_sc_hd__xor2_2
XFILLER_127_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19909_ rbzero.pov.ready_buffer\[63\] _03438_ _03558_ _03573_ vssd1 vssd1 vccd1 vccd1
+ _03574_ sky130_fd_sc_hd__a211o_1
XFILLER_102_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21802_ net328 _01391_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21733_ net259 _01322_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21664_ clknet_leaf_19_i_clk _01253_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20615_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03844_
+ sky130_fd_sc_hd__or2_1
X_21595_ clknet_leaf_70_i_clk _01184_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13920_ _07089_ _07090_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__nand2_1
X_21029_ clknet_leaf_15_i_clk _00618_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ _06959_ _06942_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__nor2_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _05382_ _05470_ _05551_ _05632_ _05958_ net37 vssd1 vssd1 vccd1 vccd1 _05979_
+ sky130_fd_sc_hd__mux4_1
XFILLER_142_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16570_ _09645_ _09659_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__xor2_1
X_13782_ _06949_ _06950_ _06952_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__nand3_1
XFILLER_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10994_ rbzero.tex_b1\[39\] rbzero.tex_b1\[40\] _04292_ vssd1 vssd1 vccd1 vccd1 _04295_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15521_ _08171_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__buf_4
X_12733_ net32 net33 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__nor2_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15452_ _08523_ _08521_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__or2b_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ rbzero.spi_registers.new_texadd\[2\]\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12664_ _05833_ net22 vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and2_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _07552_ _07573_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__xor2_1
XFILLER_208_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ _04802_ _04804_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a21oi_1
X_15383_ _08470_ _08474_ _08477_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__o21a_1
X_18171_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__nor2_1
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12595_ _03969_ gpout0.hpos\[1\] _04452_ _04628_ net16 net17 vssd1 vssd1 vccd1 vccd1
+ _05775_ sky130_fd_sc_hd__mux4_1
XFILLER_50_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17122_ _10055_ _10026_ vssd1 vssd1 vccd1 vccd1 _10142_ sky130_fd_sc_hd__or2b_1
XFILLER_204_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14334_ _07484_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11546_ rbzero.map_overlay.i_mapdy\[3\] rbzero.map_overlay.i_mapdy\[2\] rbzero.map_overlay.i_mapdy\[1\]
+ rbzero.map_overlay.i_mapdy\[0\] vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__or4_1
XFILLER_156_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17053_ _10064_ _10073_ vssd1 vssd1 vccd1 vccd1 _10074_ sky130_fd_sc_hd__xor2_1
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03791_ _03791_ vssd1 vssd1 vccd1 vccd1 clknet_0__03791_ sky130_fd_sc_hd__clkbuf_16
X_14265_ _07433_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__or2b_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11477_ rbzero.debug_overlay.playerY\[3\] vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__inv_2
XFILLER_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16004_ _09096_ _09097_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__or2_1
XFILLER_13_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13216_ _06298_ _06303_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__or2_1
X_10428_ _03995_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14196_ _07253_ _07045_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__or3_2
XFILLER_83_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20369__227 clknet_1_0__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__inv_2
XFILLER_140_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13147_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nand2_1
XFILLER_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _02212_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__xnor2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _06113_ rbzero.map_rom.i_col\[4\] _06231_ _06253_ vssd1 vssd1 vccd1 vccd1
+ _06254_ sky130_fd_sc_hd__or4b_1
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _09926_ _09927_ vssd1 vssd1 vccd1 vccd1 _09928_ sky130_fd_sc_hd__nand2_1
X_12029_ rbzero.tex_r1\[29\] _05199_ _05032_ _04890_ vssd1 vssd1 vccd1 vccd1 _05218_
+ sky130_fd_sc_hd__a31o_1
X_17886_ _02172_ _02174_ _08124_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19625_ rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\]
+ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__and4bb_1
X_16837_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09862_ sky130_fd_sc_hd__nand2_1
XFILLER_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19556_ _03406_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16768_ _09119_ _09800_ vssd1 vssd1 vccd1 vccd1 _09802_ sky130_fd_sc_hd__or2_1
XFILLER_206_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18507_ _06144_ _02724_ _09844_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
X_15719_ _08813_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__buf_4
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19487_ _03370_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16699_ rbzero.traced_texa\[-7\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a22o_1
XFILLER_179_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18438_ _02662_ _02663_ _02664_ _02665_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a211o_1
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ _05106_ _05120_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__xor2_1
XFILLER_159_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21380_ clknet_leaf_26_i_clk _00969_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22001_ net147 _01590_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20193_ _03763_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03780_ clknet_0__03780_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03780_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21716_ net242 _01305_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20474__322 clknet_1_0__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__inv_2
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21647_ clknet_leaf_82_i_clk _01236_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _03970_ _04507_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__nand2_1
X_12380_ _04937_ _05560_ _05564_ _04967_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a211o_1
XFILLER_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21578_ clknet_leaf_70_i_clk _01167_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_197_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ rbzero.spi_registers.texadd1\[15\] _04461_ _04470_ _04522_ vssd1 vssd1 vccd1
+ vccd1 _04523_ sky130_fd_sc_hd__a211o_1
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _06759_ _07219_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__or2_1
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__buf_4
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ _06175_ rbzero.wall_tracer.trackDistX\[0\] vssd1 vssd1 vccd1 vccd1 _06177_
+ sky130_fd_sc_hd__or2_1
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11193_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _04395_ vssd1 vssd1 vccd1 vccd1 _04399_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17740_ _01718_ _02029_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__or2_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _08065_ _08081_ _08082_ _08061_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__o211a_1
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13903_ _06869_ _06870_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__or2_1
XFILLER_48_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17671_ _01880_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14883_ _08032_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19410_ _04408_ _03307_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or3_2
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16622_ _09514_ _09581_ _09580_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ _07002_ _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__nand2_1
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ rbzero.color_sky\[5\] _03282_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or2_1
X_16553_ _09527_ _09537_ _09536_ vssd1 vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__a21o_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _06732_ _06792_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__nor2_1
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10977_ rbzero.tex_b1\[47\] rbzero.tex_b1\[48\] _04281_ vssd1 vssd1 vccd1 vccd1 _04286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15504_ _08513_ _08574_ _08591_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__nand3_1
X_12716_ _03969_ _04575_ _04452_ _04628_ net28 net29 vssd1 vssd1 vccd1 vccd1 _05894_
+ sky130_fd_sc_hd__mux4_1
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19272_ rbzero.spi_registers.texadd3\[5\] _03242_ vssd1 vssd1 vccd1 vccd1 _03248_
+ sky130_fd_sc_hd__or2_1
XFILLER_189_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16484_ _09554_ _09574_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__xnor2_2
X_13696_ _06799_ _06858_ _06838_ _06835_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__a22o_1
XFILLER_176_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ _02484_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15435_ _08325_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__clkinv_2
X_12647_ _05822_ _05297_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__nand2_1
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15366_ _08460_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__buf_2
X_18154_ _02424_ _02425_ _02417_ _02421_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o211a_1
X_12578_ _05729_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__nor2_2
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _10122_ _10125_ vssd1 vssd1 vccd1 vccd1 _10126_ sky130_fd_sc_hd__xor2_4
XFILLER_141_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14317_ _07486_ _07487_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__xnor2_1
X_11529_ _04707_ _04710_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and3b_1
XFILLER_184_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15297_ rbzero.wall_tracer.stepDistY\[0\] vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__inv_2
X_18085_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__or2_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17036_ _09940_ _09950_ _09949_ vssd1 vssd1 vccd1 vccd1 _10057_ sky130_fd_sc_hd__a21o_1
X_14248_ _07370_ _07416_ _07418_ _06540_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__a211o_1
XFILLER_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14179_ _07328_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__nand2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19691__69 clknet_1_0__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18987_ _02951_ _02929_ _03049_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__and3_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17938_ _02139_ _02141_ _02138_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a21bo_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17869_ _02156_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__nand2_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19608_ rbzero.spi_registers.new_texadd\[1\]\[21\] rbzero.spi_registers.spi_buffer\[21\]
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20880_ clknet_leaf_36_i_clk _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ rbzero.spi_registers.new_texadd\[0\]\[11\] rbzero.spi_registers.spi_buffer\[11\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_179_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21501_ clknet_leaf_98_i_clk _01090_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21432_ clknet_leaf_96_i_clk _01021_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21363_ clknet_leaf_22_i_clk _00952_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20317__181 clknet_1_0__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__inv_2
XFILLER_190_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21294_ clknet_leaf_33_i_clk _00883_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20176_ _03754_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ _04245_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11880_ gpout0.hpos\[6\] _04630_ _04636_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_109 vssd1 vssd1 vccd1 vccd1 ones[0] top_ew_algofoogle_109/LO sky130_fd_sc_hd__conb_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10831_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _04203_ vssd1 vssd1 vccd1 vccd1 _04209_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13550_ _06639_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__inv_2
XFILLER_186_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10762_ rbzero.tex_g1\[21\] rbzero.tex_g1\[22\] _04166_ vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12501_ _05679_ _05682_ _05640_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ _06461_ _06480_ _06603_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__mux2_1
X_10693_ _04136_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15220_ rbzero.debug_overlay.playerX\[-1\] rbzero.debug_overlay.playerX\[-2\] _08277_
+ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__or3_4
XFILLER_201_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12432_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _04913_ vssd1 vssd1 vccd1 vccd1 _05617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15151_ _08245_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__buf_2
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12363_ _05379_ _05545_ _05548_ _04650_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__a31o_1
XFILLER_154_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14102_ _07266_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__or2_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11314_ _04481_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand2_1
XFILLER_5_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15082_ rbzero.wall_tracer.stepDistY\[-3\] _08156_ _08173_ _08176_ vssd1 vssd1 vccd1
+ vccd1 _08177_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _04937_ _05475_ _05479_ _04967_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a211o_1
XFILLER_10_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _07203_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18910_ rbzero.pov.spi_buffer\[62\] rbzero.pov.ready_buffer\[62\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_101_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11245_ _04429_ _04436_ _04437_ rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 _04440_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19890_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18841_ rbzero.pov.spi_buffer\[29\] rbzero.pov.ready_buffer\[29\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _04384_ vssd1 vssd1 vccd1 vccd1 _04390_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18772_ _02961_ _02962_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__nor2_1
X_15984_ _09076_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17723_ _08428_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__nor2_1
X_14935_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.trackDistX\[1\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__mux2_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17654_ _01943_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__xnor2_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _08019_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16605_ _09561_ _09568_ _09694_ vssd1 vssd1 vccd1 vccd1 _09695_ sky130_fd_sc_hd__a21oi_1
X_13817_ _06980_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__nor2_1
X_17585_ _01803_ _01772_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__or2b_1
XFILLER_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14797_ _07826_ _07920_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__or2_1
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19324_ rbzero.floor_leak\[4\] _03272_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__or2_1
X_16536_ _09521_ _09526_ _09523_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__a21bo_1
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _06906_ _06916_ _06918_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__o21ai_2
XFILLER_17_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19255_ rbzero.spi_registers.new_texadd\[2\]\[22\] _03205_ _03236_ _03237_ vssd1
+ vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__o211a_1
X_16467_ _09556_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__xnor2_2
XFILLER_143_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__05993_ _05993_ vssd1 vssd1 vccd1 vccd1 clknet_0__05993_ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13679_ _06846_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__or2b_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _02469_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__xnor2_1
X_15418_ _08505_ _08506_ _08512_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__nand3_1
X_19186_ rbzero.spi_registers.texadd1\[17\] _03189_ vssd1 vssd1 vccd1 vccd1 _03198_
+ sky130_fd_sc_hd__or2_1
X_16398_ _09364_ _09488_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18137_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__nand2_1
XFILLER_191_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ _04464_ _06335_ _08147_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__a211o_1
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18068_ _02341_ _02350_ _02351_ _02337_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__o31a_1
XFILLER_89_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17019_ _10038_ _10039_ vssd1 vssd1 vccd1 vccd1 _10040_ sky130_fd_sc_hd__xor2_1
XFILLER_171_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20030_ _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__clkbuf_2
XFILLER_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21981_ net507 _01570_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ clknet_leaf_20_i_clk _00521_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20863_ clknet_leaf_63_i_clk _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20794_ _03968_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21415_ clknet_leaf_11_i_clk _01004_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21346_ clknet_leaf_22_i_clk _00935_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_other
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21277_ clknet_leaf_0_i_clk _00866_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11030_ _04313_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20159_ _05054_ _03737_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nand2_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12981_ _06088_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__or2_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14720_ _06568_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__or2_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11932_ _05102_ _05116_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__nor2_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _06584_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__buf_2
X_11863_ gpout0.hpos\[7\] gpout0.hpos\[8\] gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1
+ _05053_ sky130_fd_sc_hd__o21a_4
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _04121_ vssd1 vssd1 vccd1 vccd1 _04200_
+ sky130_fd_sc_hd__mux2_1
X_13602_ _06772_ _06719_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__nor2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _10327_ _10309_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__or2b_1
XFILLER_26_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _04978_ vssd1 vssd1 vccd1 vccd1 _04984_
+ sky130_fd_sc_hd__mux2_1
X_14582_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__inv_2
XFILLER_198_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16321_ _09411_ _09412_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ rbzero.tex_g1\[29\] rbzero.tex_g1\[30\] _04155_ vssd1 vssd1 vccd1 vccd1 _04164_
+ sky130_fd_sc_hd__mux2_1
X_13533_ _06474_ _06512_ _06498_ _06510_ _06589_ _06579_ vssd1 vssd1 vccd1 vccd1 _06704_
+ sky130_fd_sc_hd__mux4_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19040_ rbzero.spi_registers.new_other\[2\] _03098_ _03112_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00763_ sky130_fd_sc_hd__o211a_1
XFILLER_199_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16252_ _09126_ _09098_ _09225_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__a21oi_1
X_13464_ _06413_ _06463_ _06590_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__mux2_1
X_10676_ _04127_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12415_ _04937_ _05595_ _05599_ _04967_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a211o_1
X_15203_ _08297_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16183_ _08327_ _08384_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13395_ _06494_ _06527_ _06554_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__or4_4
XFILLER_182_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12346_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _04893_ vssd1 vssd1 vccd1 vccd1 _05532_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15134_ rbzero.wall_tracer.stepDistX\[-5\] _06261_ vssd1 vssd1 vccd1 vccd1 _08229_
+ sky130_fd_sc_hd__nor2_2
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19942_ _03436_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__and2_1
X_15065_ _08155_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__clkbuf_4
X_12277_ _04900_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__or2b_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _07133_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__nor2_1
X_11228_ _04416_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nor2_2
XFILLER_175_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19873_ _05711_ rbzero.pov.mosi_buffer\[0\] _09734_ vssd1 vssd1 vccd1 vccd1 _03549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18824_ rbzero.pov.spi_buffer\[21\] rbzero.pov.ready_buffer\[21\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02992_ sky130_fd_sc_hd__mux2_1
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _04373_ vssd1 vssd1 vccd1 vccd1 _04381_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18755_ rbzero.spi_registers.ss_buffer\[1\] _04052_ vssd1 vssd1 vccd1 vccd1 _02951_
+ sky130_fd_sc_hd__nor2_2
X_15967_ _08436_ _08479_ _09061_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__a21o_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17706_ _01939_ _01919_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__or2b_1
XFILLER_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14918_ _08036_ _08057_ _08058_ _01633_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__o211a_1
X_18686_ _09750_ _02878_ _02886_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__a21o_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _08810_ _08992_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__xnor2_2
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17637_ _08814_ _10215_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__or2_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ _06470_ _08002_ _08005_ _06516_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__a31o_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17568_ _01858_ _01859_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__and2b_1
XFILLER_189_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19307_ rbzero.spi_registers.new_texadd\[3\]\[20\] _03239_ _03267_ _03265_ vssd1
+ vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__o211a_1
XFILLER_149_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16519_ _08170_ _09608_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__or2_2
XFILLER_20_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _10059_ _09252_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19238_ rbzero.spi_registers.new_texadd\[2\]\[14\] _03221_ _03228_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__o211a_1
XFILLER_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20535__377 clknet_1_1__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__inv_2
XFILLER_165_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19169_ _03173_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21200_ clknet_leaf_21_i_clk _00789_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21131_ clknet_leaf_96_i_clk _00720_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21062_ clknet_leaf_82_i_clk _00651_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20013_ rbzero.pov.ready_buffer\[58\] _03586_ _03617_ _03652_ vssd1 vssd1 vccd1 vccd1
+ _03653_ sky130_fd_sc_hd__o211a_1
XFILLER_8_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20429__282 clknet_1_0__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__inv_2
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21964_ net490 _01553_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20280__147 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__inv_2
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ clknet_leaf_69_i_clk _00504_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21895_ net421 _01484_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ clknet_leaf_56_i_clk _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03462_ clknet_0__03462_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03462_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20777_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__or2_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ rbzero.tex_r1\[1\] rbzero.tex_r1\[2\] _04046_ vssd1 vssd1 vccd1 vccd1 _04049_
+ sky130_fd_sc_hd__mux2_1
XFILLER_210_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ _04012_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12200_ rbzero.tex_g1\[12\] _04906_ _05181_ _05385_ _05386_ vssd1 vssd1 vccd1 vccd1
+ _05387_ sky130_fd_sc_hd__a311o_1
XFILLER_182_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ rbzero.wall_tracer.visualWallDist\[-2\] _06327_ _04443_ vssd1 vssd1 vccd1
+ vccd1 _06351_ sky130_fd_sc_hd__a21o_1
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12131_ _04903_ _05304_ _05309_ _05318_ _04887_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__o311a_1
X_21329_ clknet_leaf_33_i_clk _00918_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ rbzero.tex_r1\[57\] _05199_ _05182_ _04952_ vssd1 vssd1 vccd1 vccd1 _05251_
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ rbzero.tex_b1\[30\] rbzero.tex_b1\[31\] _04303_ vssd1 vssd1 vccd1 vccd1 _04305_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _09641_ _09611_ vssd1 vssd1 vccd1 vccd1 _09892_ sky130_fd_sc_hd__or2b_1
XFILLER_78_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _08827_ _08915_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__nor2_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _02746_ _02750_ _02751_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _08250_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__clkbuf_4
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12964_ rbzero.wall_tracer.visualWallDist\[-1\] rbzero.wall_tracer.visualWallDist\[-2\]
+ rbzero.wall_tracer.visualWallDist\[-3\] _06139_ vssd1 vssd1 vccd1 vccd1 _06140_
+ sky130_fd_sc_hd__or4_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14703_ _07872_ _07858_ _07806_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ rbzero.wall_tracer.rayAddendX\[9\] _02527_ _09760_ _02693_ _02696_ vssd1
+ vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__o221a_1
X_11915_ _05099_ _05101_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or3_1
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15683_ _08776_ _08777_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__or2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _06020_ _06048_ _05999_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__a21o_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _01694_ _01714_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ _07529_ _07802_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__xnor2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ rbzero.row_render.texu\[0\] _05034_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_
+ sky130_fd_sc_hd__or3b_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _10369_ _10371_ vssd1 vssd1 vccd1 vccd1 _10372_ sky130_fd_sc_hd__nand2_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04889_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__buf_6
X_14565_ _07698_ _07726_ _07731_ _07733_ _07735_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__a32oi_4
XFILLER_158_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16304_ _09394_ _09395_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10728_ _04143_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__clkbuf_4
X_13516_ _06469_ _06683_ _06684_ _06686_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__o2bb2a_4
X_17284_ _10301_ _10302_ vssd1 vssd1 vccd1 vccd1 _10303_ sky130_fd_sc_hd__nor2_1
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _07645_ _07665_ _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__a21boi_1
X_19023_ _03084_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__clkbuf_4
X_16235_ _09326_ _09327_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__05761_ _05761_ vssd1 vssd1 vccd1 vccd1 clknet_0__05761_ sky130_fd_sc_hd__clkbuf_16
X_10659_ _04118_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13447_ _06494_ _06527_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__nor2_1
XFILLER_103_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16166_ _09257_ _09258_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__nand2_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _06463_ _06518_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nor2_1
XFILLER_115_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ _08162_ _08206_ _08211_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__o21ai_2
XFILLER_177_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _05009_ vssd1 vssd1 vccd1 vccd1 _05515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _08145_ _09187_ _09189_ _09190_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__o31ai_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19925_ _03116_ _03556_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__nor2_1
X_15048_ _08142_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19856_ _03540_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18807_ rbzero.pov.spi_buffer\[13\] rbzero.pov.ready_buffer\[13\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02983_ sky130_fd_sc_hd__mux2_1
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19787_ _03504_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16999_ _09907_ _09909_ _09906_ vssd1 vssd1 vccd1 vccd1 _10020_ sky130_fd_sc_hd__o21ba_1
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18738_ _02474_ _02475_ _02476_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a31oi_2
XFILLER_110_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18669_ _02794_ _05132_ _02868_ _02869_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__nor4_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20700_ _03913_ _03914_ _03915_ _03908_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a22o_1
X_21680_ clknet_leaf_0_i_clk _01269_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20631_ _03854_ _03855_ _03856_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a21o_1
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19712__87 clknet_1_0__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21114_ clknet_leaf_94_i_clk _00703_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21045_ clknet_leaf_86_i_clk _00634_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21947_ net473 _01536_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11700_ _04814_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__buf_4
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05841_ _05844_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__o21ba_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21878_ net404 _01467_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11631_ _04820_ _04794_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nor2_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ clknet_leaf_50_i_clk _00418_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11562_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] _04751_ vssd1
+ vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a21o_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14350_ _07446_ _07478_ _07497_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__a31o_1
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10513_ rbzero.tex_r1\[9\] rbzero.tex_r1\[10\] _04035_ vssd1 vssd1 vccd1 vccd1 _04040_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13301_ _06386_ _06391_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__nor2_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14281_ _07446_ _07451_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__or2_1
X_11493_ _04666_ _04669_ _04678_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__and4b_1
XFILLER_13_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13232_ rbzero.wall_tracer.visualWallDist\[-1\] _06327_ _04443_ vssd1 vssd1 vccd1
+ vccd1 _06403_ sky130_fd_sc_hd__a21oi_1
X_16020_ _09105_ _09106_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__and2_1
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10444_ rbzero.tex_r1\[42\] rbzero.tex_r1\[43\] _04002_ vssd1 vssd1 vccd1 vccd1 _04004_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13163_ _06321_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _05010_ vssd1 vssd1 vccd1 vccd1 _05302_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17971_ _02258_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__inv_2
X_13094_ _06267_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19710_ clknet_1_1__leaf__04634_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__buf_1
XFILLER_123_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16922_ _09941_ _09942_ _09943_ vssd1 vssd1 vccd1 vccd1 _09944_ sky130_fd_sc_hd__a21o_1
X_12045_ rbzero.tex_r1\[38\] _05031_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or2_1
XFILLER_46_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20219__92 clknet_1_1__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
X_19641_ rbzero.pov.spi_counter\[6\] _03454_ _03446_ vssd1 vssd1 vccd1 vccd1 _03456_
+ sky130_fd_sc_hd__a21boi_1
X_16853_ _09874_ _09875_ _09876_ vssd1 vssd1 vccd1 vccd1 _09877_ sky130_fd_sc_hd__and3_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _08835_ _08858_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_0__f__05879_ clknet_0__05879_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05879_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19572_ _03414_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
X_16784_ _06105_ _09810_ _09811_ _09812_ _09815_ vssd1 vssd1 vccd1 vccd1 _09816_ sky130_fd_sc_hd__o311a_1
XFILLER_19_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13996_ _07130_ _07142_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__nor2_1
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18523_ rbzero.debug_overlay.playerX\[4\] _02736_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02737_ sky130_fd_sc_hd__mux2_1
X_15735_ _08815_ _08829_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__nor2_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12947_ rbzero.debug_overlay.playerX\[2\] _06120_ _06121_ rbzero.debug_overlay.playerY\[4\]
+ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a221o_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _02569_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__inv_2
X_15666_ _08758_ _08760_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__nor2_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _06028_ _06018_ _06024_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__and3_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _01697_ _10288_ _08476_ _09044_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__or4_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07746_ _07787_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__nor2_2
X_11829_ rbzero.row_render.wall\[1\] rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1
+ vccd1 _05019_ sky130_fd_sc_hd__or2b_1
X_18385_ _05106_ _05120_ _02614_ _02615_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15597_ _08685_ _08691_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _10352_ _10354_ vssd1 vssd1 vccd1 vccd1 _10355_ sky130_fd_sc_hd__nor2_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14548_ _07675_ _07718_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__nand2_1
XFILLER_202_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17267_ _10284_ _10285_ vssd1 vssd1 vccd1 vccd1 _10286_ sky130_fd_sc_hd__xor2_1
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14479_ _07252_ _07361_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__nor2_1
XFILLER_88_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19006_ _03088_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__clkbuf_1
X_16218_ rbzero.wall_tracer.visualWallDist\[-11\] _08149_ _09310_ vssd1 vssd1 vccd1
+ vccd1 _09311_ sky130_fd_sc_hd__and3_1
XFILLER_128_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ _10204_ _10217_ vssd1 vssd1 vccd1 vccd1 _10218_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ rbzero.wall_tracer.visualWallDist\[7\] _08475_ vssd1 vssd1 vccd1 vccd1 _09242_
+ sky130_fd_sc_hd__nand2_4
XFILLER_103_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20311__176 clknet_1_1__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__inv_2
X_19908_ _08239_ _03570_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__nor2_1
XFILLER_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19839_ _03531_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21801_ net327 _01390_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21732_ net258 _01321_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21663_ clknet_leaf_19_i_clk _01252_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20614_ rbzero.texV\[-5\] _03814_ _03819_ _03843_ vssd1 vssd1 vccd1 vccd1 _01606_
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21594_ clknet_leaf_69_i_clk _01183_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20392__248 clknet_1_1__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__inv_2
XFILLER_165_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20545_ clknet_1_0__leaf__04634_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__buf_1
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19697__75 clknet_1_1__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
XFILLER_165_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20286__153 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__inv_2
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21028_ clknet_leaf_16_i_clk _00617_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _07019_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12801_ _05958_ _05297_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nand2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ _04294_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
X_13781_ _06757_ _06738_ _06951_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__and3_1
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15520_ _08611_ _08604_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__or2b_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12732_ _05899_ _05881_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__nor2_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15451_ _08534_ _08536_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__o21ai_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__nor2_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14402_ _07554_ _07571_ _07572_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18170_ _01868_ _02439_ _02364_ rbzero.wall_tracer.trackDistY\[5\] vssd1 vssd1 vccd1
+ vccd1 _00566_ sky130_fd_sc_hd__o2bb2a_1
X_11614_ _04746_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15382_ _08476_ _08461_ _08459_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__or3b_1
XFILLER_184_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _04589_ _04704_ _04419_ _03973_ _05763_ net17 vssd1 vssd1 vccd1 vccd1 _05774_
+ sky130_fd_sc_hd__mux4_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _10029_ _10054_ vssd1 vssd1 vccd1 vccd1 _10141_ sky130_fd_sc_hd__nand2_1
XFILLER_196_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20451__301 clknet_1_1__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__inv_2
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14333_ _07252_ _07249_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__nor2_1
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11545_ _04652_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__inv_2
XFILLER_204_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17052_ _10071_ _10072_ vssd1 vssd1 vccd1 vccd1 _10073_ sky130_fd_sc_hd__and2b_1
XFILLER_156_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03790_ _03790_ vssd1 vssd1 vccd1 vccd1 clknet_0__03790_ sky130_fd_sc_hd__clkbuf_16
XFILLER_167_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14264_ _07432_ _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__xnor2_1
X_11476_ _04662_ _04663_ _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a22o_1
XFILLER_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_88_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16003_ _09096_ _09097_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__nand2_1
X_10427_ rbzero.tex_r1\[50\] rbzero.tex_r1\[51\] _03991_ vssd1 vssd1 vccd1 vccd1 _03995_
+ sky130_fd_sc_hd__mux2_1
X_13215_ _06379_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__or2_1
XFILLER_100_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _07302_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__clkbuf_2
XFILLER_139_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13146_ _06310_ _06312_ _06316_ _06285_ _06286_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__o2111ai_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17954_ _02213_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__xnor2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ rbzero.map_rom.f1 rbzero.map_rom.c6 rbzero.map_rom.a6 _06121_ vssd1 vssd1
+ vccd1 vccd1 _06253_ sky130_fd_sc_hd__and4_1
X_16905_ _09898_ _09899_ _09925_ vssd1 vssd1 vccd1 vccd1 _09927_ sky130_fd_sc_hd__nand3_1
X_12028_ rbzero.tex_r1\[31\] _05195_ _05216_ _04923_ vssd1 vssd1 vccd1 vccd1 _05217_
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17885_ _01972_ _01980_ _02077_ _02078_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a31o_1
XFILLER_38_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16836_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09861_ sky130_fd_sc_hd__nor2_1
X_19624_ rbzero.pov.spi_counter\[5\] rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\]
+ rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__and4bb_1
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19555_ rbzero.spi_registers.new_texadd\[0\]\[19\] rbzero.spi_registers.spi_buffer\[19\]
+ _03380_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16767_ _09119_ _09800_ vssd1 vssd1 vccd1 vccd1 _09801_ sky130_fd_sc_hd__nand2_1
XFILLER_94_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13979_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__inv_2
XFILLER_111_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18506_ rbzero.debug_overlay.playerX\[0\] _06108_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02724_ sky130_fd_sc_hd__mux2_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15718_ _08328_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19486_ rbzero.spi_registers.new_mapd\[7\] rbzero.spi_registers.spi_buffer\[7\] _03362_
+ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__mux2_1
XFILLER_202_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16698_ rbzero.traced_texa\[-8\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] rbzero.wall_tracer.rayAddendX\[4\]
+ rbzero.wall_tracer.rayAddendX\[3\] _02597_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__o41a_1
XFILLER_179_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _08722_ _08717_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18368_ _02582_ _02586_ _02599_ _02600_ _08136_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a311oi_1
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17319_ _10332_ _10337_ vssd1 vssd1 vccd1 vccd1 _10338_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18299_ rbzero.wall_tracer.rayAddendX\[-4\] _02527_ _02533_ _02537_ vssd1 vssd1 vccd1
+ vccd1 _00597_ sky130_fd_sc_hd__o22a_1
XFILLER_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22000_ net146 _01589_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
X_20192_ rbzero.spi_registers.new_texadd\[3\]\[11\] rbzero.spi_registers.spi_buffer\[11\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__mux2_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21715_ net241 _01304_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21646_ clknet_leaf_80_i_clk _01235_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21577_ clknet_leaf_94_i_clk _01166_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11330_ rbzero.spi_registers.texadd3\[15\] _04465_ _04456_ rbzero.spi_registers.texadd2\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a22o_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11261_ _03969_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__inv_2
XFILLER_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13000_ _06175_ rbzero.wall_tracer.trackDistX\[0\] _06173_ rbzero.wall_tracer.trackDistX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__a22o_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11192_ _04398_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14951_ rbzero.wall_tracer.visualWallDist\[6\] _08046_ vssd1 vssd1 vccd1 vccd1 _08082_
+ sky130_fd_sc_hd__or2_1
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13902_ _07071_ _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__xnor2_2
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17670_ _01958_ _01960_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__xor2_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14882_ rbzero.wall_tracer.stepDistY\[10\] _08031_ _07868_ vssd1 vssd1 vccd1 vccd1
+ _08032_ sky130_fd_sc_hd__mux2_1
X_16621_ _09642_ _09710_ vssd1 vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13833_ _06955_ _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__and2_1
XFILLER_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ rbzero.color_sky\[4\] _03280_ _03286_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__a21o_1
X_16552_ _09611_ _09641_ vssd1 vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__xnor2_1
X_13764_ _06790_ _06733_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__nor2_1
X_10976_ _04285_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _08593_ _08597_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__xnor2_1
X_12715_ _04589_ _04704_ _04419_ _03973_ _05881_ _05888_ vssd1 vssd1 vccd1 vccd1 _05893_
+ sky130_fd_sc_hd__mux4_1
X_19271_ rbzero.spi_registers.new_texadd\[3\]\[4\] _03240_ _03247_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00859_ sky130_fd_sc_hd__o211a_1
XFILLER_206_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16483_ _09572_ _09573_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__xor2_2
XFILLER_203_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ _06820_ _06822_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__nand2_1
XFILLER_188_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18222_ rbzero.spi_registers.new_texadd\[2\]\[2\] _02483_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15434_ _08250_ _08251_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__and2b_1
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ _05824_ net26 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__nor2_1
XFILLER_180_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18153_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nor2_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ rbzero.wall_tracer.visualWallDist\[-11\] _08156_ vssd1 vssd1 vccd1 vccd1
+ _08460_ sky130_fd_sc_hd__nand2_1
XFILLER_129_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ net15 _05752_ _05713_ _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a22o_2
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ _10123_ _10009_ _10124_ vssd1 vssd1 vccd1 vccd1 _10125_ sky130_fd_sc_hd__o21ai_2
XFILLER_184_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _07433_ _07435_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__xnor2_1
X_18084_ _09837_ _02365_ _02340_ rbzero.wall_tracer.trackDistY\[-7\] vssd1 vssd1 vccd1
+ vccd1 _00554_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11528_ _04711_ _04712_ _04715_ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__and4_1
XFILLER_184_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15296_ rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__inv_2
XFILLER_8_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17035_ _10026_ _10055_ vssd1 vssd1 vccd1 vccd1 _10056_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19676__56 clknet_1_1__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
X_14247_ _07417_ _07398_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__nor2_1
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11459_ _04646_ _04647_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__o21a_1
XFILLER_125_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14178_ _07311_ _07330_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__o21ai_1
XFILLER_139_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__xnor2_4
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _03077_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__clkbuf_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__xnor2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17868_ _02120_ _02155_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__or2_1
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ _03432_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16819_ _06184_ _09786_ _09846_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a21oi_1
X_17799_ _02025_ _02086_ _02087_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a21o_1
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20458__307 clknet_1_1__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__inv_2
X_19538_ _03397_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19469_ rbzero.spi_registers.spi_cmd\[0\] _02474_ _03974_ _03350_ vssd1 vssd1 vccd1
+ vccd1 _03360_ sky130_fd_sc_hd__and4b_1
XFILLER_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21500_ clknet_leaf_98_i_clk _01089_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21431_ clknet_leaf_96_i_clk _01020_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21362_ clknet_leaf_21_i_clk _00951_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21293_ clknet_leaf_33_i_clk _00882_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20175_ rbzero.spi_registers.new_texadd\[3\]\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__mux2_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _04208_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20398__254 clknet_1_0__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__inv_2
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10761_ _04172_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12500_ _05680_ _05681_ _05661_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__mux2_1
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10692_ rbzero.tex_g1\[54\] rbzero.tex_g1\[55\] _04132_ vssd1 vssd1 vccd1 vccd1 _04136_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13480_ _06618_ _06536_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__nand2_1
XFILLER_205_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12431_ _04919_ _05611_ _05615_ _04889_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a211o_1
XFILLER_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21629_ clknet_leaf_88_i_clk _01218_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15150_ _06262_ _08240_ _08244_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__o21ai_4
X_12362_ _04702_ _04743_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__or3_1
XFILLER_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ _07227_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ rbzero.texu_hot\[4\] _04480_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__or2_1
X_12293_ _05476_ _05477_ _05478_ _05190_ _04952_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__o221a_1
X_15081_ _08160_ _08175_ vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__nor2_1
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14032_ _07161_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__xnor2_1
X_11244_ _04436_ _04437_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__and3_1
XFILLER_153_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11175_ _04389_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__clkbuf_1
X_18840_ _02967_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18771_ rbzero.spi_registers.spi_counter\[5\] _02959_ _02951_ vssd1 vssd1 vccd1 vccd1
+ _02962_ sky130_fd_sc_hd__o21ai_1
X_15983_ _08619_ _09077_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__nor2_1
XFILLER_121_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17722_ rbzero.wall_tracer.visualWallDist\[6\] _08421_ vssd1 vssd1 vccd1 vccd1 _02012_
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14934_ _08065_ _08068_ _08070_ _08061_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__o211a_1
XFILLER_209_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17653_ _09542_ _01718_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__nor2_1
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ rbzero.wall_tracer.stepDistY\[6\] _08018_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08019_ sky130_fd_sc_hd__mux2_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _09562_ _09567_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__nor2_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13816_ _06979_ _06975_ _06978_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__and3_1
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17584_ _01872_ _01873_ _09866_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a21o_1
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14796_ _07822_ _07879_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__and2_1
XFILLER_32_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ rbzero.spi_registers.new_leak\[3\] _03271_ _03276_ _03265_ vssd1 vssd1 vccd1
+ vccd1 _00882_ sky130_fd_sc_hd__o211a_1
X_16535_ _09498_ _09501_ _09624_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__a21bo_1
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13747_ _06777_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
X_10959_ _04276_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19254_ _03212_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__clkbuf_4
X_16466_ _08434_ _09186_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__nor2_1
XFILLER_148_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _06846_ _06847_ _06848_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__or3_1
X_18205_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__xor2_1
X_15417_ _08510_ _08511_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12629_ net47 _05801_ _05790_ _05780_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__o211a_1
X_19185_ rbzero.spi_registers.new_texadd\[1\]\[16\] _03188_ _03196_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__o211a_1
X_16397_ _09008_ _09242_ vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__nor2_1
XFILLER_185_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18136_ _10011_ _02410_ _02340_ rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1
+ vccd1 _00561_ sky130_fd_sc_hd__o2bb2a_1
X_15348_ _04464_ _06037_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__nor2_1
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18067_ _02348_ _02349_ _02347_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21a_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15279_ _08235_ _08373_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__nor2_1
XFILLER_171_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17018_ _09008_ _09890_ vssd1 vssd1 vccd1 vccd1 _10039_ sky130_fd_sc_hd__nand2_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ rbzero.spi_registers.spi_buffer\[15\] rbzero.spi_registers.spi_buffer\[14\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ net506 _01569_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20931_ clknet_leaf_54_i_clk _00520_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20862_ clknet_leaf_61_i_clk _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20793_ _03110_ _03966_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__and3_1
XFILLER_168_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21414_ clknet_leaf_1_i_clk _01003_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21345_ clknet_leaf_9_i_clk _00934_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21276_ clknet_leaf_1_i_clk _00865_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20158_ _04670_ _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nand2_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20089_ _05106_ _03676_ _03698_ _03695_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a211o_1
X_12980_ rbzero.map_overlay.i_mapdy\[0\] _06130_ _06089_ rbzero.map_overlay.i_mapdy\[1\]
+ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__o221a_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ rbzero.debug_overlay.vplaneX\[-6\] vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20406__261 clknet_1_0__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__inv_2
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14650_ _07818_ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__nand2_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _04661_ _05049_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__o21ai_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _06771_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__clkbuf_4
X_10813_ _04199_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14581_ _07749_ _07751_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__xor2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04979_ _04980_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_14_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16320_ _08373_ _08497_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__nor2_1
X_13532_ _06598_ _06607_ _06614_ _06647_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a22oi_4
X_10744_ _04163_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _09342_ _09343_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__and2_2
XFILLER_186_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13463_ _06574_ _06628_ _06630_ _06631_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__a2111o_1
XFILLER_201_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10675_ rbzero.tex_g1\[62\] rbzero.tex_g1\[63\] _04046_ vssd1 vssd1 vccd1 vccd1 _04127_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15202_ _08292_ _08162_ _08296_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__a21o_1
XFILLER_199_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12414_ _04944_ _05596_ _05598_ _04919_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o211a_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16182_ _09273_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13394_ _06545_ _06558_ _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__nor3_2
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__buf_2
XFILLER_154_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12345_ _04826_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__or2_1
XFILLER_127_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19941_ rbzero.debug_overlay.playerX\[3\] _03594_ vssd1 vssd1 vccd1 vccd1 _03598_
+ sky130_fd_sc_hd__or2_1
X_15064_ _07892_ _08144_ _08154_ _08158_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__o211a_2
X_12276_ rbzero.color_sky\[3\] rbzero.color_floor\[3\] _04825_ vssd1 vssd1 vccd1 vccd1
+ _05463_ sky130_fd_sc_hd__mux2_1
XFILLER_107_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14015_ _07132_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__xor2_1
X_11227_ _04421_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19872_ _03548_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18823_ _02991_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
X_11158_ _04380_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15966_ _08469_ _08478_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__nor2_1
X_11089_ _04344_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__clkbuf_1
X_18754_ _02943_ _02944_ _02946_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__and4_1
XFILLER_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17705_ _01893_ _01913_ _01911_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a21o_1
X_14917_ rbzero.wall_tracer.visualWallDist\[-4\] _08047_ vssd1 vssd1 vccd1 vccd1 _08058_
+ sky130_fd_sc_hd__or2_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ _08809_ _08866_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__nor2_1
X_18685_ rbzero.wall_tracer.rayAddendY\[6\] _09751_ _02885_ _08136_ vssd1 vssd1 vccd1
+ vccd1 _02886_ sky130_fd_sc_hd__a22o_1
XFILLER_48_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17636_ _01925_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__and2_1
XFILLER_64_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14848_ _07826_ _08003_ _08004_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__a21o_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _01856_ _01857_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__nand2_1
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ rbzero.wall_tracer.stepDistY\[-6\] _07944_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07945_ sky130_fd_sc_hd__mux2_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16518_ rbzero.wall_tracer.visualWallDist\[10\] _08475_ vssd1 vssd1 vccd1 vccd1 _09608_
+ sky130_fd_sc_hd__nand2_1
X_19306_ rbzero.spi_registers.texadd3\[20\] _03241_ vssd1 vssd1 vccd1 vccd1 _03267_
+ sky130_fd_sc_hd__or2_1
XFILLER_143_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _01788_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__nand2_1
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16449_ _09518_ _09539_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__xor2_1
X_19237_ rbzero.spi_registers.texadd2\[14\] _03222_ vssd1 vssd1 vccd1 vccd1 _03228_
+ sky130_fd_sc_hd__or2_1
XFILLER_158_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19168_ rbzero.spi_registers.new_texadd\[1\]\[9\] _03174_ _03187_ _03184_ vssd1 vssd1
+ vccd1 vccd1 _00816_ sky130_fd_sc_hd__o211a_1
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20234__106 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__inv_2
XFILLER_9_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18119_ _02386_ _02389_ _02387_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__o21ai_1
X_19099_ rbzero.spi_registers.new_texadd\[0\]\[3\] _03141_ _03148_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00786_ sky130_fd_sc_hd__o211a_1
XFILLER_172_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03808_ _03808_ vssd1 vssd1 vccd1 vccd1 clknet_0__03808_ sky130_fd_sc_hd__clkbuf_16
X_21130_ clknet_leaf_93_i_clk _00719_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21061_ clknet_leaf_98_i_clk _00650_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20012_ _06114_ _03648_ _03437_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__a21o_1
XFILLER_98_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21963_ net489 _01552_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20914_ clknet_leaf_69_i_clk _00503_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21894_ net420 _01483_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ clknet_leaf_66_i_clk _00434_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_0__f__03461_ clknet_0__03461_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03461_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20776_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__nand2_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ rbzero.tex_r1\[34\] rbzero.tex_r1\[35\] _04002_ vssd1 vssd1 vccd1 vccd1 _04012_
+ sky130_fd_sc_hd__mux2_1
XFILLER_149_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20436__287 clknet_1_0__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__inv_2
X_10391_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__buf_4
XFILLER_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _04941_ _05312_ _05317_ _04955_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a211o_1
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21328_ clknet_leaf_30_i_clk _00917_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ rbzero.tex_r1\[59\] _05002_ _05249_ _04922_ vssd1 vssd1 vccd1 vccd1 _05250_
+ sky130_fd_sc_hd__o211a_1
X_21259_ clknet_leaf_100_i_clk _00848_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _04304_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15820_ _08910_ _08344_ _08911_ _08914_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__o31a_1
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15751_ _08276_ _08440_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__nor2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ rbzero.wall_tracer.visualWallDist\[3\] rbzero.wall_tracer.visualWallDist\[2\]
+ rbzero.wall_tracer.visualWallDist\[1\] rbzero.wall_tracer.visualWallDist\[0\] vssd1
+ vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__or4_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14702_ _07850_ _07852_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _02682_ _02685_ _02695_ _04434_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a211o_1
X_11914_ _05093_ _05102_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__nor2_1
X_15682_ _08771_ _08772_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12894_ _06044_ _06045_ _06053_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__a211o_1
XFILLER_79_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17421_ _01696_ _01713_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__xor2_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _07471_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__xnor2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ rbzero.row_render.texu\[4\] rbzero.row_render.texu\[3\] _05024_ _04889_ vssd1
+ vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__a31o_1
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _10370_ vssd1 vssd1 vccd1 vccd1 _10371_ sky130_fd_sc_hd__inv_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14564_ _07734_ _07731_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__xnor2_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11776_ _04912_ _04962_ _04963_ _04965_ _04940_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__o221a_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16303_ _08368_ _08535_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__or2_1
XFILLER_53_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ _06641_ _06606_ _06685_ _06669_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__a211oi_2
XFILLER_207_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17283_ _10299_ _10300_ vssd1 vssd1 vccd1 vccd1 _10302_ sky130_fd_sc_hd__and2_1
X_10727_ _04154_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__clkbuf_1
X_14495_ _07646_ _07664_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__or2b_1
XFILLER_174_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19022_ rbzero.map_overlay.i_otherx\[0\] _03101_ vssd1 vssd1 vccd1 vccd1 _03102_
+ sky130_fd_sc_hd__or2_1
X_16234_ _09323_ _09325_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__and2_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ _06581_ _06596_ _06601_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__o211ai_4
X_10658_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _04110_ vssd1 vssd1 vccd1 vccd1 _04118_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16165_ _09256_ _09254_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__or2b_1
XFILLER_186_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13377_ _06546_ _06547_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__nand2_1
X_10589_ rbzero.tex_r0\[40\] rbzero.tex_r0\[39\] _04077_ vssd1 vssd1 vccd1 vccd1 _04082_
+ sky130_fd_sc_hd__mux2_1
XFILLER_103_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15116_ rbzero.debug_overlay.playerX\[-7\] _08185_ _08210_ _06261_ vssd1 vssd1 vccd1
+ vccd1 _08211_ sky130_fd_sc_hd__a211o_1
X_12328_ _04953_ _05509_ _05513_ _04967_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a211o_1
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ _08144_ _08452_ _08453_ _08405_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__a31oi_4
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19924_ rbzero.debug_overlay.playerX\[-1\] _03559_ _03583_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01175_ sky130_fd_sc_hd__a211o_1
X_15047_ _04430_ _08141_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__nor2_1
X_12259_ rbzero.tex_g1\[38\] _04830_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19855_ rbzero.pov.spi_buffer\[64\] rbzero.pov.spi_buffer\[65\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18806_ _02982_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19786_ rbzero.pov.spi_buffer\[31\] rbzero.pov.spi_buffer\[32\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XFILLER_209_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16998_ _09928_ _09897_ vssd1 vssd1 vccd1 vccd1 _10019_ sky130_fd_sc_hd__or2b_1
XFILLER_37_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18737_ _02475_ rbzero.spi_registers.spi_cmd\[3\] _02932_ vssd1 vssd1 vccd1 vccd1
+ _02933_ sky130_fd_sc_hd__and3b_1
X_15949_ _09043_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18668_ _02794_ _05132_ _02868_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__o22a_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ _01785_ _01793_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18599_ _02802_ _02805_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__xor2_1
XFILLER_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20630_ _03854_ _03855_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nand3_1
XFILLER_177_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21113_ clknet_leaf_94_i_clk _00702_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21044_ clknet_leaf_86_i_clk _00633_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21946_ net472 _01535_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21877_ net403 _01466_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _04760_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__inv_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20828_ clknet_leaf_50_i_clk _00417_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11561_ rbzero.texV\[8\] _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__and3_1
X_20518__362 clknet_1_1__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__inv_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20759_ rbzero.wall_tracer.rayAddendX\[-7\] _02606_ _02557_ _03946_ vssd1 vssd1 vccd1
+ vccd1 _01649_ sky130_fd_sc_hd__a22o_1
XFILLER_204_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13300_ _06365_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__clkinv_2
X_10512_ _04039_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__clkbuf_1
X_14280_ _07447_ _07450_ _06540_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11492_ _04679_ _04628_ _04419_ _04680_ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__o221a_1
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _06394_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_2
X_10443_ _04003_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13162_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__nand2_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _04933_ vssd1 vssd1 vccd1 vccd1 _05301_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17970_ _02256_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nor2_1
X_13093_ rbzero.wall_tracer.mapY\[6\] _06078_ _06101_ vssd1 vssd1 vccd1 vccd1 _06268_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_105_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16921_ _08327_ _09176_ _09037_ _08813_ vssd1 vssd1 vccd1 vccd1 _09943_ sky130_fd_sc_hd__o22a_1
XFILLER_151_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ rbzero.tex_r1\[40\] _04935_ _05195_ _05231_ _05232_ vssd1 vssd1 vccd1 vccd1
+ _05233_ sky130_fd_sc_hd__a311o_1
XFILLER_104_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19640_ _03454_ _03455_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__nor2_1
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16852_ _09861_ _09864_ _09862_ vssd1 vssd1 vccd1 vccd1 _09876_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15803_ _08896_ _08897_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__nand2_1
X_16783_ _08123_ _09813_ _09814_ vssd1 vssd1 vccd1 vccd1 _09815_ sky130_fd_sc_hd__or3_1
X_19571_ rbzero.spi_registers.new_texadd\[1\]\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
X_20263__132 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__inv_2
XFILLER_20_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ _07112_ _07143_ _07165_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__a21oi_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15734_ _08816_ _08344_ _08826_ _08827_ _08828_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__o41a_1
X_18522_ _09775_ _09774_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__xnor2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ rbzero.debug_overlay.playerX\[3\] rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1
+ _06122_ sky130_fd_sc_hd__xor2_1
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15665_ _08708_ _08709_ _08759_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__o21a_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18453_ _02678_ _02679_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__nor2_1
XFILLER_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12877_ _06048_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and2_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ rbzero.wall_tracer.visualWallDist\[1\] _08421_ vssd1 vssd1 vccd1 vccd1 _01697_
+ sky130_fd_sc_hd__nand2_2
X_14616_ _07741_ _07747_ _07748_ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__or4b_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _04957_ _04977_ _04996_ _05016_ _05017_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o221a_2
X_18384_ _05106_ _05120_ _02614_ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__and4bb_1
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15596_ _08689_ _08690_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__nand2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _10201_ _10227_ _10353_ vssd1 vssd1 vccd1 vccd1 _10354_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14547_ _07253_ _07444_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__nor2_1
X_11759_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _04948_ vssd1 vssd1 vccd1 vccd1 _04949_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266_ _09005_ _09687_ vssd1 vssd1 vccd1 vccd1 _10285_ sky130_fd_sc_hd__and2_1
XFILLER_186_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14478_ _07606_ _07613_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19005_ net46 rbzero.spi_registers.sclk_buffer\[0\] _09734_ vssd1 vssd1 vccd1 vccd1
+ _03088_ sky130_fd_sc_hd__mux2_1
X_16217_ _08145_ _09308_ _09309_ _09190_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__o31a_2
XFILLER_162_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13429_ _06544_ _06499_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__nand2_4
X_17197_ _09970_ _09972_ _08431_ vssd1 vssd1 vccd1 vccd1 _10217_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ _09162_ _09240_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__nand2_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _09171_ _09172_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19907_ rbzero.debug_overlay.playerX\[-6\] _03569_ _03572_ _03302_ vssd1 vssd1 vccd1
+ vccd1 _01170_ sky130_fd_sc_hd__o211a_1
XFILLER_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19838_ rbzero.pov.spi_buffer\[56\] rbzero.pov.spi_buffer\[57\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 i_debug_map_overlay vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
X_19769_ rbzero.pov.spi_buffer\[23\] rbzero.pov.spi_buffer\[24\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XFILLER_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21800_ net326 _01389_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21731_ net257 _01320_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21662_ clknet_leaf_19_i_clk _01251_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20613_ _03840_ _03842_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__xnor2_1
X_21593_ clknet_leaf_69_i_clk _01182_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21027_ clknet_leaf_16_i_clk _00616_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_43_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ _05952_ net38 vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__nor2_1
XFILLER_74_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13780_ _06790_ _06755_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__nor2_1
X_10992_ rbzero.tex_b1\[40\] rbzero.tex_b1\[41\] _04292_ vssd1 vssd1 vccd1 vccd1 _04294_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12731_ net31 net30 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nor2_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21929_ net455 _01518_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _08543_ _08544_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__nand2_1
X_12662_ _05824_ _05829_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__nand2_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14401_ _07555_ _07570_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__nor2_1
XFILLER_204_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11613_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _04803_
+ sky130_fd_sc_hd__xor2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15381_ _08475_ _08445_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__nand2_1
X_12593_ _05770_ _05766_ _05772_ net20 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17120_ _10138_ _10139_ vssd1 vssd1 vccd1 vccd1 _10140_ sky130_fd_sc_hd__nand2_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14332_ _07501_ _07502_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11544_ _04670_ rbzero.map_overlay.i_mapdy\[4\] rbzero.map_overlay.i_mapdy\[2\] _04731_
+ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a22oi_1
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17051_ _10068_ _10070_ vssd1 vssd1 vccd1 vccd1 _10072_ sky130_fd_sc_hd__nand2_1
XFILLER_13_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14263_ _06993_ _07248_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nor2_1
XFILLER_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ _04652_ rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 _04665_
+ sky130_fd_sc_hd__or2_1
X_16002_ _08659_ _08761_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__and2_1
XFILLER_13_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13214_ rbzero.wall_tracer.rcp_sel\[0\] _06382_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_
+ sky130_fd_sc_hd__a21oi_4
X_10426_ _03994_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14194_ _07342_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__inv_2
XFILLER_3_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17953_ _02215_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__xnor2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ rbzero.map_rom.f1 rbzero.map_rom.c6 rbzero.map_rom.a6 rbzero.map_rom.f2 _06251_
+ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__a221o_1
X_16904_ _09898_ _09899_ _09925_ vssd1 vssd1 vccd1 vccd1 _09926_ sky130_fd_sc_hd__a21o_1
X_12027_ rbzero.tex_r1\[30\] _05182_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__or2_1
X_17884_ _01972_ _01980_ _02077_ _02078_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a311o_1
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19623_ rbzero.pov.spi_counter\[0\] _03439_ rbzero.pov.spi_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 _03443_ sky130_fd_sc_hd__a21o_1
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16835_ _06182_ _09785_ _09860_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19554_ _03405_ vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _07101_ _07103_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__nor2_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16766_ rbzero.wall_tracer.mapX\[10\] _09799_ vssd1 vssd1 vccd1 vccd1 _09800_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _02723_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
X_15717_ _08782_ _08806_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__buf_6
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19485_ _03369_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
X_16697_ rbzero.traced_texa\[-9\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__a22o_1
XFILLER_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _02637_ _02638_ _02650_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__nor3_1
X_15648_ _08678_ _08729_ _08742_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__nand3_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15579_ _08195_ _08201_ _08234_ _08213_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__o22ai_1
X_18367_ _02582_ _02586_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17318_ _10335_ _10336_ vssd1 vssd1 vccd1 vccd1 _10337_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _02534_ _02535_ _02536_ _09745_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a31o_1
XFILLER_30_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17249_ _10157_ _10158_ _10155_ _10156_ vssd1 vssd1 vccd1 vccd1 _10268_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20191_ _03762_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ net240 _01303_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20400__256 clknet_1_0__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__inv_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ clknet_leaf_80_i_clk _01234_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_36_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21576_ clknet_leaf_95_i_clk _01165_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11260_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__buf_4
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11191_ rbzero.tex_b0\[10\] rbzero.tex_b0\[9\] _04395_ vssd1 vssd1 vccd1 vccd1 _04398_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20481__328 clknet_1_1__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__inv_2
X_14950_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.trackDistX\[6\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__mux2_1
XFILLER_47_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22059_ clknet_leaf_79_i_clk _01648_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13901_ _06807_ _06861_ _06852_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14881_ _07891_ _06541_ _06631_ _07998_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__and4bb_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16620_ _09708_ _09709_ vssd1 vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__and2b_1
X_13832_ _06953_ _06954_ _06947_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__a21o_1
XFILLER_210_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16551_ _09639_ _09640_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__nand2_1
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13763_ _06893_ _06892_ _06891_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__a21o_1
X_10975_ rbzero.tex_b1\[48\] rbzero.tex_b1\[49\] _04281_ vssd1 vssd1 vccd1 vccd1 _04285_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15502_ _08594_ _08596_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__xor2_1
X_12714_ _05889_ _05885_ _05891_ net32 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a22o_1
X_16482_ _09436_ _09438_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__and2_1
X_19270_ rbzero.spi_registers.texadd3\[4\] _03242_ vssd1 vssd1 vccd1 vccd1 _03247_
+ sky130_fd_sc_hd__or2_1
X_13694_ _06862_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__xor2_2
XFILLER_44_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15433_ _08495_ _08527_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18221_ rbzero.spi_registers.spi_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__buf_4
X_12645_ net25 vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__inv_2
XFILLER_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20375__233 clknet_1_1__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__inv_2
XFILLER_203_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15364_ _08455_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__nor2_2
XFILLER_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18152_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__and2_1
XFILLER_168_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12576_ _05726_ _05754_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a21o_2
XFILLER_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17103_ _09717_ _10005_ vssd1 vssd1 vccd1 vccd1 _10124_ sky130_fd_sc_hd__nand2_1
X_14315_ _07252_ _07249_ _07484_ _07485_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__o31ai_2
XFILLER_157_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18083_ _09872_ _02363_ _02364_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__o21a_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11527_ rbzero.map_overlay.i_otherx\[3\] _04410_ _04411_ _04705_ _04716_ vssd1 vssd1
+ vccd1 vccd1 _04717_ sky130_fd_sc_hd__o221a_1
X_15295_ _08195_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17034_ _10029_ _10054_ vssd1 vssd1 vccd1 vccd1 _10055_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _06785_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _03985_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14177_ _07308_ _07329_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__or2_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11389_ _04458_ _04521_ _04524_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__or3_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nand2_2
XFILLER_140_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ rbzero.spi_registers.spi_buffer\[23\] rbzero.spi_registers.spi_buffer\[22\]
+ _03051_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17936_ _10059_ _09890_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__nand2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ rbzero.map_overlay.i_othery\[0\] _06130_ vssd1 vssd1 vccd1 vccd1 _06235_
+ sky130_fd_sc_hd__nor2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17867_ _02120_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__nand2_1
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19606_ rbzero.spi_registers.new_texadd\[1\]\[20\] rbzero.spi_registers.spi_buffer\[20\]
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
X_16818_ _09842_ _09843_ _09844_ _09845_ vssd1 vssd1 vccd1 vccd1 _09846_ sky130_fd_sc_hd__o211a_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _02003_ _02004_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19537_ rbzero.spi_registers.new_texadd\[0\]\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16749_ _09783_ vssd1 vssd1 vccd1 vccd1 _09786_ sky130_fd_sc_hd__clkbuf_4
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ rbzero.spi_registers.got_new_vinf _03118_ _03316_ _03358_ vssd1 vssd1 vccd1
+ vccd1 _00944_ sky130_fd_sc_hd__a31o_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ rbzero.wall_tracer.rayAddendX\[5\] _09745_ _02648_ _02534_ vssd1 vssd1 vccd1
+ vccd1 _02649_ sky130_fd_sc_hd__a22o_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19399_ _02483_ rbzero.spi_registers.new_floor\[2\] _03319_ vssd1 vssd1 vccd1 vccd1
+ _03322_ sky130_fd_sc_hd__mux2_1
XFILLER_50_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21430_ clknet_leaf_96_i_clk _01019_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21361_ clknet_leaf_21_i_clk _00950_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20312_ clknet_1_1__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__buf_1
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21292_ clknet_leaf_31_i_clk _00881_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20174_ _03753_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_72_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_87_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ rbzero.tex_g1\[22\] rbzero.tex_g1\[23\] _04166_ vssd1 vssd1 vccd1 vccd1 _04172_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10691_ _04135_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12430_ _04827_ _05612_ _05613_ _05614_ _04939_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o221a_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21628_ clknet_leaf_88_i_clk _01217_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12361_ _05546_ _05290_ _05465_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__o21a_1
XFILLER_193_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21559_ clknet_leaf_90_i_clk _01148_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14100_ _07226_ _07267_ _07268_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__or4bb_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _04501_ _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__or2_1
X_15080_ _04463_ _06053_ _08142_ _08174_ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_25_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12292_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _05009_ vssd1 vssd1 vccd1 vccd1 _05478_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14031_ _07162_ _07201_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__xor2_2
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11243_ rbzero.trace_state\[3\] _04429_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_175_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ rbzero.tex_b0\[18\] rbzero.tex_b0\[17\] _04384_ vssd1 vssd1 vccd1 vccd1 _04389_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19681__60 clknet_1_1__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18770_ rbzero.spi_registers.spi_counter\[5\] _02959_ vssd1 vssd1 vccd1 vccd1 _02961_
+ sky130_fd_sc_hd__and2_1
X_15982_ _08164_ _09076_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__or2_1
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17721_ _02008_ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__nand2_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14933_ _08069_ _08035_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__nand2_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _01942_ _10093_ _01832_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__or3b_1
XFILLER_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14864_ _06470_ _06575_ _07874_ _08017_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__a31o_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _09686_ _09692_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13815_ _06981_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17583_ _01872_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__nor2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14795_ _07822_ _07886_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__nor2_1
XFILLER_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19322_ rbzero.floor_leak\[3\] _03272_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or2_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16534_ _09371_ _09499_ vssd1 vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__nand2_1
X_13746_ _06790_ _06769_ _06719_ _06772_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__o22a_1
X_10958_ rbzero.tex_b1\[56\] rbzero.tex_b1\[57\] _04270_ vssd1 vssd1 vccd1 vccd1 _04276_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19253_ rbzero.spi_registers.texadd2\[22\] _03207_ vssd1 vssd1 vccd1 vccd1 _03236_
+ sky130_fd_sc_hd__or2_1
X_16465_ _09545_ _09555_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__xnor2_1
X_13677_ _06766_ _06781_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__xnor2_1
X_10889_ rbzero.tex_g0\[26\] rbzero.tex_g0\[25\] _04237_ vssd1 vssd1 vccd1 vccd1 _04240_
+ sky130_fd_sc_hd__mux2_1
XFILLER_177_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18204_ _02455_ _02464_ _02465_ _02462_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a31o_1
XFILLER_188_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15416_ _08368_ _08228_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__nor2_1
X_12628_ _05792_ _05804_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__nor2_1
X_16396_ _09244_ _09364_ vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__nand2_1
X_19184_ _03110_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18135_ _02341_ _02408_ _02409_ _02339_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__o31a_1
X_15347_ _08000_ _08425_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__xor2_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12559_ _04651_ _04657_ _05652_ _05653_ net10 net12 vssd1 vssd1 vccd1 vccd1 _05740_
+ sky130_fd_sc_hd__mux4_1
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15278_ _08287_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18066_ _02347_ _02348_ _02349_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__nor3_1
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17017_ _10035_ _10037_ vssd1 vssd1 vccd1 vccd1 _10038_ sky130_fd_sc_hd__xnor2_1
X_14229_ _07329_ _07399_ _07332_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__o21ai_1
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _03068_ vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _01840_ _02093_ _02205_ _02206_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__o22a_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18899_ rbzero.pov.spi_buffer\[57\] rbzero.pov.ready_buffer\[57\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_113_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20930_ clknet_leaf_54_i_clk _00519_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20861_ clknet_leaf_65_i_clk _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20792_ gpout4.clk_div\[0\] gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__or2_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21413_ clknet_leaf_12_i_clk _01002_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21344_ clknet_leaf_9_i_clk _00933_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21275_ clknet_leaf_7_i_clk _00864_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20157_ _05645_ _03739_ _03742_ _03118_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__o211a_1
XFILLER_77_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ rbzero.pov.ready_buffer\[18\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__and3_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ rbzero.debug_overlay.vplaneX\[-8\] _05117_ _05118_ rbzero.debug_overlay.vplaneX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a22o_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ rbzero.trace_state\[0\] _05050_ _04635_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a21o_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06633_ _06650_ _06654_ _06655_ _06657_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__a32oi_4
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ rbzero.tex_g0\[62\] rbzero.tex_g0\[61\] _04121_ vssd1 vssd1 vccd1 vccd1 _04199_
+ sky130_fd_sc_hd__mux2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _07727_ _07750_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__xor2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11792_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__buf_4
XFILLER_25_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _06619_ _06676_ _06602_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__o21ai_2
X_10743_ rbzero.tex_g1\[30\] rbzero.tex_g1\[31\] _04155_ vssd1 vssd1 vccd1 vccd1 _04163_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _09222_ _09224_ _09340_ _09341_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _06632_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__buf_4
XFILLER_201_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _04126_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ rbzero.wall_tracer.stepDistY\[-8\] _08157_ _08293_ _08295_ vssd1 vssd1 vccd1
+ vccd1 _08296_ sky130_fd_sc_hd__a2bb2o_4
X_12413_ _04981_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__or2_1
X_16181_ _09005_ _08553_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__nor2_1
XFILLER_166_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13393_ _06370_ _06544_ _06559_ _06521_ _06563_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__a41o_1
XFILLER_194_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _06262_ _08219_ _08226_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__o21ai_4
X_12344_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _04907_ vssd1 vssd1 vccd1 vccd1 _05530_
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19940_ rbzero.debug_overlay.playerX\[2\] _03569_ _03597_ _03579_ vssd1 vssd1 vccd1
+ vccd1 _01178_ sky130_fd_sc_hd__o211a_1
X_15063_ _08157_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__buf_4
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20487__334 clknet_1_1__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__inv_2
XFILLER_154_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ _05457_ _05461_ _04900_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__or3b_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ _06733_ _06719_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__or2_1
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _04412_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand2_1
XFILLER_175_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19871_ rbzero.pov.spi_buffer\[72\] rbzero.pov.spi_buffer\[73\] _03467_ vssd1 vssd1
+ vccd1 vccd1 _03548_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18822_ rbzero.pov.spi_buffer\[20\] rbzero.pov.ready_buffer\[20\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02991_ sky130_fd_sc_hd__mux2_1
X_11157_ rbzero.tex_b0\[26\] rbzero.tex_b0\[25\] _04373_ vssd1 vssd1 vccd1 vccd1 _04380_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18753_ rbzero.spi_registers.spi_counter\[3\] _02948_ vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__xnor2_1
X_15965_ _09041_ _09059_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__xnor2_2
X_11088_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _04340_ vssd1 vssd1 vccd1 vccd1 _04344_
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17704_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__nor2_1
XFILLER_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14916_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.trackDistX\[-4\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__mux2_1
X_18684_ _02883_ _02884_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _08865_ _08903_ _08905_ _08990_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__a22o_2
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _09662_ _01922_ _01924_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14847_ _06574_ _07977_ _07978_ _06631_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__a31o_1
XFILLER_17_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _01856_ _01857_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__nor2_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14778_ _07891_ _07942_ _07943_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__or3_2
XFILLER_147_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19305_ rbzero.spi_registers.new_texadd\[3\]\[19\] _03254_ _03266_ _03265_ vssd1
+ vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__o211a_1
XFILLER_210_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16517_ _09605_ _09606_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__nor2_1
X_13729_ _06889_ _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__and2b_1
XFILLER_56_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17497_ _10315_ _09079_ _01787_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__o21ai_1
XFILLER_177_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19236_ rbzero.spi_registers.new_texadd\[2\]\[13\] _03221_ _03227_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__o211a_1
X_16448_ _09527_ _09538_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19167_ rbzero.spi_registers.texadd1\[9\] _03176_ vssd1 vssd1 vccd1 vccd1 _03187_
+ sky130_fd_sc_hd__or2_1
X_16379_ _09467_ _09469_ vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__and2_1
XFILLER_30_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18118_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__nand2_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19098_ rbzero.spi_registers.texadd0\[3\] _03143_ vssd1 vssd1 vccd1 vccd1 _03148_
+ sky130_fd_sc_hd__or2_1
XFILLER_117_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03807_ _03807_ vssd1 vssd1 vccd1 vccd1 clknet_0__03807_ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18049_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__nor2_1
XFILLER_105_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21060_ clknet_leaf_98_i_clk _00649_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20011_ _06114_ _03649_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nor2_1
XFILLER_141_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19660__41 clknet_1_0__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21962_ net488 _01551_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20913_ clknet_leaf_69_i_clk _00502_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21893_ net419 _01482_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20844_ clknet_leaf_66_i_clk _00433_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03460_ clknet_0__03460_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03460_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20775_ gpout1.clk_div\[0\] net63 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nor2_1
XFILLER_167_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__buf_4
XFILLER_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21327_ clknet_leaf_30_i_clk _00916_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ rbzero.tex_r1\[58\] _05031_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or2_1
XFILLER_46_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21258_ clknet_leaf_0_i_clk _00847_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ rbzero.tex_b1\[31\] rbzero.tex_b1\[32\] _04303_ vssd1 vssd1 vccd1 vccd1 _04304_
+ sky130_fd_sc_hd__mux2_1
X_20209_ _03771_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21189_ clknet_leaf_22_i_clk _00778_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _08529_ _08733_ _08844_ _08790_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__a22o_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12962_ rbzero.wall_tracer.visualWallDist\[7\] rbzero.wall_tracer.visualWallDist\[6\]
+ rbzero.wall_tracer.visualWallDist\[5\] rbzero.wall_tracer.visualWallDist\[4\] vssd1
+ vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__or4_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _04411_ _05080_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__or2_1
X_14701_ _07806_ _07850_ _07853_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__and3_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _08287_ _08358_ _08774_ _08775_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__o31a_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12893_ _06055_ _06056_ _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__or3_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _01711_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__nand2_1
XFILLER_61_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ rbzero.row_render.texu\[4\] rbzero.row_render.texu\[3\] _05022_ _04889_ vssd1
+ vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__o31a_1
X_14632_ _07530_ _07802_ _07527_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__o21ba_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _10265_ _10242_ _10368_ vssd1 vssd1 vccd1 vccd1 _10370_ sky130_fd_sc_hd__and3_1
XFILLER_202_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14563_ _07698_ _07726_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__nand2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ rbzero.tex_r0\[26\] _04964_ _04934_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a21o_1
XFILLER_53_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16302_ _09276_ _09393_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__xnor2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10726_ rbzero.tex_g1\[38\] rbzero.tex_g1\[39\] _04144_ vssd1 vssd1 vccd1 vccd1 _04154_
+ sky130_fd_sc_hd__mux2_1
X_13514_ _06576_ _06659_ _06660_ _06619_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__o211a_1
X_17282_ _10299_ _10300_ vssd1 vssd1 vccd1 vccd1 _10301_ sky130_fd_sc_hd__nor2_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14494_ _07646_ _07664_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19021_ rbzero.spi_registers.got_new_other _03100_ vssd1 vssd1 vccd1 vccd1 _03101_
+ sky130_fd_sc_hd__and2_2
X_16233_ _09323_ _09325_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__nor2_1
X_13445_ _06602_ _06611_ _06615_ _06469_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__a211o_1
X_10657_ _04117_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _09254_ _09256_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__or2b_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _06442_ _06444_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__and2_1
X_10588_ _04081_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ _05190_ _05510_ _05511_ _05512_ _04890_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__o221a_1
X_15115_ _08185_ _08209_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__nor2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16095_ _08012_ _08450_ _09188_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__nor3_1
XFILLER_182_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19923_ _04409_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__clkbuf_4
X_15046_ rbzero.trace_state\[3\] rbzero.trace_state\[2\] vssd1 vssd1 vccd1 vccd1 _08141_
+ sky130_fd_sc_hd__nand2_1
X_12258_ rbzero.tex_g1\[40\] _04905_ _04910_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1
+ _05445_ sky130_fd_sc_hd__a311o_1
XFILLER_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11209_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _04054_ vssd1 vssd1 vccd1 vccd1 _04407_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19854_ _03539_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
X_12189_ rbzero.color_sky\[2\] rbzero.color_floor\[2\] _04825_ vssd1 vssd1 vccd1 vccd1
+ _05377_ sky130_fd_sc_hd__mux2_1
XFILLER_1_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18805_ rbzero.pov.spi_buffer\[12\] rbzero.pov.ready_buffer\[12\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19785_ _03503_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
X_16997_ _10017_ _10003_ vssd1 vssd1 vccd1 vccd1 _10018_ sky130_fd_sc_hd__nand2_2
XFILLER_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18736_ rbzero.spi_registers.spi_cmd\[0\] _02474_ vssd1 vssd1 vccd1 vccd1 _02932_
+ sky130_fd_sc_hd__nand2_1
XFILLER_114_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15948_ _08455_ _09042_ _08357_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__a21o_1
XFILLER_3_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20541__383 clknet_1_0__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__inv_2
XFILLER_37_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18667_ _02821_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _02869_
+ sky130_fd_sc_hd__and2_1
X_15879_ _08960_ _08962_ _08966_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__o21a_1
XFILLER_184_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20240__111 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__inv_2
X_17618_ _01792_ _01786_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__and2b_1
XFILLER_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18598_ _02803_ _02804_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__nand2_1
XFILLER_205_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17549_ _01839_ _01840_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__and2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19219_ rbzero.spi_registers.new_texadd\[2\]\[6\] _03206_ _03217_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00837_ sky130_fd_sc_hd__o211a_1
XFILLER_177_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11444__1 clknet_1_1__leaf__04634_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
XFILLER_30_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21112_ clknet_leaf_94_i_clk _00701_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21043_ clknet_leaf_86_i_clk _00632_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_141_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21945_ net471 _01534_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ net402 _01465_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ clknet_leaf_50_i_clk _00416_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11560_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _04750_ sky130_fd_sc_hd__or2_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20758_ _02517_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ rbzero.tex_r1\[10\] rbzero.tex_r1\[11\] _04035_ vssd1 vssd1 vccd1 vccd1 _04039_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11491_ rbzero.debug_overlay.playerX\[4\] _03972_ vssd1 vssd1 vccd1 vccd1 _04681_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20689_ _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__xnor2_1
XFILLER_137_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13230_ _06310_ _06312_ _06316_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or3_1
X_10442_ rbzero.tex_r1\[43\] rbzero.tex_r1\[44\] _04002_ vssd1 vssd1 vccd1 vccd1 _04003_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _06324_ _06328_ _06331_ _06322_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a31oi_4
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _04650_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__inv_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ rbzero.wall_tracer.mapY\[7\] _06077_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__xor2_1
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16920_ _08327_ _09037_ vssd1 vssd1 vccd1 vccd1 _09942_ sky130_fd_sc_hd__nor2_1
X_12043_ rbzero.tex_r1\[41\] _05199_ _05032_ _04952_ vssd1 vssd1 vccd1 vccd1 _05232_
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16851_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09875_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15802_ _08870_ _08894_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__xor2_1
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19570_ _03413_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_1
X_16782_ _08905_ _08990_ vssd1 vssd1 vccd1 vccd1 _09814_ sky130_fd_sc_hd__nor2_1
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13994_ _07144_ _07110_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__and2b_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18521_ _02735_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
X_15733_ _08821_ _08825_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__or2b_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__inv_2
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _02662_ _02667_ _02677_ _08135_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a31o_1
X_15664_ _08661_ _08707_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__or2_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _06049_ _06050_ _06007_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__a211o_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _10332_ _10337_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a21bo_1
XFILLER_18_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14615_ _07723_ _07737_ _07783_ _07784_ _07785_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__a221oi_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ net42 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__clkinv_4
X_18383_ rbzero.debug_overlay.vplaneX\[-1\] _05111_ vssd1 vssd1 vccd1 vccd1 _02615_
+ sky130_fd_sc_hd__nand2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15595_ _08673_ _08686_ _08688_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__nand3_1
X_20552__13 clknet_1_0__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
XFILLER_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _10224_ _10226_ vssd1 vssd1 vccd1 vccd1 _10353_ sky130_fd_sc_hd__and2b_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11758_ _04908_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__clkbuf_8
X_14546_ _07685_ _07705_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10709_ _04145_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__clkbuf_1
X_17265_ _10282_ _10283_ vssd1 vssd1 vccd1 vccd1 _10284_ sky130_fd_sc_hd__xor2_1
XFILLER_146_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14477_ _07638_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__xnor2_1
X_11689_ _04866_ _04877_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21oi_1
X_19004_ _03087_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__clkbuf_1
X_16216_ _08012_ _08450_ _09188_ _08023_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__o31a_1
X_13428_ _06495_ _06578_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__nor2_2
X_17196_ _09167_ _10215_ vssd1 vssd1 vccd1 vccd1 _10216_ sky130_fd_sc_hd__nor2_1
XFILLER_128_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16147_ _09164_ _09144_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__or2b_1
XFILLER_154_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ _06507_ _06466_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__or3_1
XFILLER_182_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _08373_ _08384_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__nor2_1
XFILLER_29_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19906_ rbzero.pov.ready_buffer\[62\] _03438_ _03559_ _03571_ vssd1 vssd1 vccd1 vccd1
+ _03572_ sky130_fd_sc_hd__a211o_1
X_15029_ _06159_ _06233_ _08126_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__or3_1
XFILLER_142_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19837_ _03530_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19768_ _03494_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
Xinput2 i_debug_trace_overlay vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20225__97 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__inv_2
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18719_ _02894_ _02903_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nor2_1
X_19699_ clknet_1_0__leaf__03457_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__buf_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21730_ net256 _01319_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21661_ clknet_leaf_19_i_clk _01250_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20612_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _03841_ vssd1 vssd1 vccd1 vccd1
+ _03842_ sky130_fd_sc_hd__o21ai_1
XFILLER_123_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21592_ clknet_leaf_15_i_clk _01181_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21026_ clknet_leaf_15_i_clk _00615_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_2
XFILLER_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20247__117 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__inv_2
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991_ _04293_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ net51 net41 net40 _05263_ _05888_ _05881_ vssd1 vssd1 vccd1 vccd1 _05908_
+ sky130_fd_sc_hd__mux4_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21928_ net454 _01517_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _05833_ _05834_ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a21oi_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21859_ net385 _01448_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _04748_ _04752_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__a21o_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _07555_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__xor2_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15380_ _08149_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__buf_4
X_12592_ net17 _05770_ net19 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14331_ _07426_ _07425_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__or2b_1
X_11543_ _04648_ _04730_ rbzero.map_overlay.i_mapdy\[2\] _04731_ _04732_ vssd1 vssd1
+ vccd1 vccd1 _04733_ sky130_fd_sc_hd__o221a_1
X_20293__159 clknet_1_0__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__inv_2
XFILLER_183_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17050_ _10068_ _10070_ vssd1 vssd1 vccd1 vccd1 _10071_ sky130_fd_sc_hd__nor2_1
XFILLER_52_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14262_ _07316_ _07209_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__or2_1
XFILLER_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11474_ _04653_ rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 _04664_
+ sky130_fd_sc_hd__nand2_1
X_16001_ _09093_ _09095_ vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__xor2_1
X_13213_ _04427_ _06063_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ rbzero.tex_r1\[51\] rbzero.tex_r1\[52\] _03991_ vssd1 vssd1 vccd1 vccd1 _03994_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14193_ _07211_ _07251_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__or2_1
XFILLER_139_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13144_ _06313_ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nand2_1
XFILLER_152_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _02225_ _02239_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__xnor2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13075_ _06228_ _06089_ _06107_ _06120_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__a221o_1
XFILLER_183_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16903_ _09910_ _09924_ vssd1 vssd1 vccd1 vccd1 _09925_ sky130_fd_sc_hd__xnor2_1
X_12026_ rbzero.tex_r1\[16\] _04906_ _05181_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1
+ _05215_ sky130_fd_sc_hd__a311o_1
X_17883_ _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__inv_2
X_19622_ rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\] _03439_ vssd1 vssd1
+ vccd1 vccd1 _03442_ sky130_fd_sc_hd__and3_1
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16834_ _06105_ _09857_ _09858_ _09812_ _09859_ vssd1 vssd1 vccd1 vccd1 _09860_ sky130_fd_sc_hd__o311a_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19553_ rbzero.spi_registers.new_texadd\[0\]\[18\] rbzero.spi_registers.spi_buffer\[18\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
X_16765_ rbzero.wall_tracer.mapX\[9\] _09119_ _09798_ vssd1 vssd1 vccd1 vccd1 _09799_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13977_ _07145_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18504_ rbzero.wall_tracer.mapY\[5\] _02722_ _02704_ vssd1 vssd1 vccd1 vccd1 _02723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15716_ _08809_ _08810_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__nand2_1
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19484_ rbzero.spi_registers.new_mapd\[6\] rbzero.spi_registers.spi_buffer\[6\] _03362_
+ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__mux2_1
X_12928_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__buf_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16696_ _09753_ vssd1 vssd1 vccd1 vccd1 _09756_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18435_ _02597_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _02663_
+ sky130_fd_sc_hd__or2_1
XFILLER_206_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15647_ _08738_ _08741_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__nand2_1
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12859_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18366_ _02598_ rbzero.wall_tracer.rayAddendX\[2\] vssd1 vssd1 vccd1 vccd1 _02599_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_187_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15578_ _08212_ _08201_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__or3_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17317_ _09406_ _09677_ vssd1 vssd1 vccd1 vccd1 _10336_ sky130_fd_sc_hd__nor2_1
X_14529_ _07690_ _07691_ _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__a21o_1
X_18297_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__or2_1
XFILLER_147_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20352__212 clknet_1_1__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__inv_2
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _10178_ _10147_ vssd1 vssd1 vccd1 vccd1 _10267_ sky130_fd_sc_hd__or2b_1
XFILLER_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ _10188_ _10198_ vssd1 vssd1 vccd1 vccd1 _10199_ sky130_fd_sc_hd__xor2_1
XFILLER_162_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20190_ rbzero.spi_registers.new_texadd\[3\]\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__mux2_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21713_ net239 _01302_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21644_ clknet_leaf_80_i_clk _01233_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21575_ clknet_leaf_95_i_clk _01164_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_40 _06217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20457_ clknet_1_1__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__buf_1
XFILLER_118_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ _04397_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22058_ clknet_leaf_79_i_clk _01647_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21009_ clknet_leaf_78_i_clk _00598_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13900_ _07069_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xor2_2
XFILLER_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14880_ _08030_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_i_clk clknet_1_1_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13831_ _06992_ _07001_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__or2b_1
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16550_ _09612_ _09613_ _09638_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__nand3_1
X_10974_ _04284_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
X_13762_ _06893_ _06891_ _06892_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__nand3_1
XFILLER_44_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15501_ _08595_ _08518_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__xor2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12713_ _05888_ _05889_ net31 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a21oi_1
X_16481_ _09558_ _09571_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13693_ _06834_ _06839_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a21bo_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _02482_ vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__clkbuf_1
X_15432_ _08515_ _08525_ _08526_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__a21o_1
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12644_ _05822_ _05057_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__or2_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18151_ _10259_ _02423_ _02364_ rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1
+ vccd1 _00563_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_169_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15363_ _08457_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__buf_4
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12575_ gpout1.clk_div\[1\] _05749_ _05755_ clknet_1_0__leaf__04634_ _05721_ vssd1
+ vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__o221a_2
XFILLER_180_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17102_ _09717_ _10005_ vssd1 vssd1 vccd1 vccd1 _10123_ sky130_fd_sc_hd__nor2_1
XFILLER_184_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14314_ _07482_ _07483_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__nand2_1
XFILLER_200_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18082_ _02336_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ rbzero.map_overlay.i_otherx\[0\] _04412_ vssd1 vssd1 vccd1 vccd1 _04716_
+ sky130_fd_sc_hd__xnor2_1
X_15294_ _08387_ _08388_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _10040_ _10053_ vssd1 vssd1 vccd1 vccd1 _10054_ sky130_fd_sc_hd__xor2_1
X_14245_ _07344_ _07369_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__or2_1
X_11457_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _04647_ sky130_fd_sc_hd__or3_2
XFILLER_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10408_ rbzero.tex_r1\[59\] rbzero.tex_r1\[60\] _03980_ vssd1 vssd1 vccd1 vccd1 _03985_
+ sky130_fd_sc_hd__mux2_1
X_14176_ _07345_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__nand2_1
XFILLER_139_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11388_ _04419_ _04568_ _04577_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a31o_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13127_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nor2_1
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _03076_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17935_ _02221_ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__xnor2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ rbzero.map_overlay.i_otherx\[4\] vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__inv_2
XFILLER_140_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12009_ _04817_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__buf_4
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17866_ _02121_ _02154_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16817_ _09822_ _09101_ vssd1 vssd1 vccd1 vccd1 _09845_ sky130_fd_sc_hd__nand2_1
X_19605_ _03431_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__clkbuf_1
X_17797_ _02027_ _01995_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__or2b_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19536_ _03396_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16748_ _09779_ _09780_ _09784_ _09785_ rbzero.wall_tracer.mapX\[6\] vssd1 vssd1
+ vccd1 vccd1 _00523_ sky130_fd_sc_hd__a32o_1
XFILLER_35_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19467_ _03359_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16679_ rbzero.row_render.size\[6\] _09746_ _09750_ _07975_ vssd1 vssd1 vccd1 vccd1
+ _00489_ sky130_fd_sc_hd__a22o_1
XFILLER_146_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18418_ _02646_ _02647_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19398_ _03321_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18349_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__or2_1
XFILLER_148_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21360_ clknet_leaf_22_i_clk _00949_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667__47 clknet_1_0__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
X_21291_ clknet_leaf_33_i_clk _00880_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20173_ rbzero.spi_registers.new_texadd\[3\]\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__mux2_1
XFILLER_107_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20359__218 clknet_1_0__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__inv_2
XFILLER_197_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ rbzero.tex_g1\[55\] rbzero.tex_g1\[56\] _04132_ vssd1 vssd1 vccd1 vccd1 _04135_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21627_ clknet_leaf_88_i_clk _01216_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ _05277_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__inv_2
XFILLER_139_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21558_ clknet_leaf_70_i_clk _01147_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _04485_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__nand2_1
XFILLER_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12291_ rbzero.tex_b0\[62\] _04978_ _05198_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a21o_1
X_21489_ net207 _01078_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _07199_ _07200_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__and2_1
X_11242_ rbzero.trace_state\[0\] vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__buf_2
XFILLER_175_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11173_ _04388_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15981_ rbzero.wall_tracer.visualWallDist\[5\] _08149_ vssd1 vssd1 vccd1 vccd1 _09076_
+ sky130_fd_sc_hd__nand2_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ rbzero.wall_tracer.visualWallDist\[5\] _01699_ _02009_ vssd1 vssd1 vccd1
+ vccd1 _02010_ sky130_fd_sc_hd__a21o_1
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14932_ rbzero.wall_tracer.visualWallDist\[0\] vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__inv_2
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _08889_ _08816_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__and2_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14863_ _07989_ _07889_ _06516_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__a21o_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _06433_ _09687_ _09691_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__mux2_1
X_13814_ _06754_ _06983_ _06984_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17582_ _01761_ _01763_ _01762_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__o21ba_1
XFILLER_21_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14794_ _07903_ _07956_ _07957_ _07941_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__a211o_1
XFILLER_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19321_ rbzero.spi_registers.new_leak\[2\] _03271_ _03275_ _03265_ vssd1 vssd1 vccd1
+ vccd1 _00881_ sky130_fd_sc_hd__o211a_1
XFILLER_204_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16533_ _09620_ _09622_ vssd1 vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__xor2_1
X_13745_ _06901_ _06903_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__a211oi_1
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10957_ _04275_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20299__165 clknet_1_1__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__inv_2
XFILLER_182_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19252_ rbzero.spi_registers.new_texadd\[2\]\[21\] _03205_ _03235_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__o211a_1
XFILLER_71_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16464_ _09195_ _09421_ _08431_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__a21oi_1
X_13676_ _06845_ _06844_ _06819_ _06816_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__a211oi_1
X_10888_ _04239_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
X_18203_ _02262_ _02468_ _02364_ rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1
+ vccd1 _00570_ sky130_fd_sc_hd__o2bb2a_1
X_15415_ _08508_ _08509_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__nand2_1
XFILLER_129_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ net55 _05791_ _05802_ net53 _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a221o_1
X_19183_ rbzero.spi_registers.texadd1\[16\] _03189_ vssd1 vssd1 vccd1 vccd1 _03196_
+ sky130_fd_sc_hd__or2_1
X_16395_ _09404_ _09385_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__or2b_1
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18134_ _02401_ _02403_ _02406_ _02407_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__o211a_1
XFILLER_89_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15346_ _08440_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _05731_ _05736_ _05738_ _05717_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__o31a_1
XFILLER_185_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18065_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__and2_1
XFILLER_8_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11509_ gpout0.hpos\[6\] gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or2_1
X_15277_ _08368_ _08369_ _08371_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12489_ net43 _05637_ _05638_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a31o_1
XFILLER_176_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17016_ _09008_ _09491_ _09901_ _10036_ vssd1 vssd1 vccd1 vccd1 _10037_ sky130_fd_sc_hd__o31a_1
XFILLER_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14228_ _07306_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nor2_1
XFILLER_160_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14159_ _07308_ _07329_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__nand2_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20464__313 clknet_1_0__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__inv_2
XFILLER_140_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ rbzero.spi_registers.spi_buffer\[14\] rbzero.spi_registers.spi_buffer\[13\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17918_ _10221_ _01729_ _02093_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__and3_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18898_ _03030_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17849_ _02009_ _02137_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__nand2_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20860_ clknet_leaf_62_i_clk _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ _03387_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__clkbuf_1
X_20791_ gpout4.clk_div\[0\] gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__nand2_1
XFILLER_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21412_ clknet_leaf_2_i_clk _01001_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21343_ clknet_leaf_9_i_clk _00932_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21274_ clknet_leaf_7_i_clk _00863_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20330__192 clknet_1_1__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__inv_2
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20156_ _05645_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nand2_1
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20087_ rbzero.pov.ready_buffer\[17\] _03684_ _03697_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01225_ sky130_fd_sc_hd__o211a_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ rbzero.trace_state\[3\] _04429_ _04436_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and3_4
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _04198_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__clkbuf_1
X_11791_ _04817_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__buf_4
XFILLER_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20989_ clknet_leaf_25_i_clk _00578_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ _06641_ _06672_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__nor2_1
X_10742_ _04162_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ rbzero.tex_g1\[63\] net50 _04046_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__mux2_1
X_13461_ _06448_ _06467_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__nand2_4
XFILLER_185_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15200_ _08143_ _08294_ _08160_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__a21oi_1
X_12412_ rbzero.tex_b1\[15\] rbzero.tex_b1\[14\] _04913_ vssd1 vssd1 vccd1 vccd1 _05597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16180_ _09271_ _09272_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__nand2_1
XFILLER_166_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _06448_ _06467_ _06483_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__and4_1
XFILLER_138_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15131_ rbzero.wall_tracer.visualWallDist\[-6\] _08158_ _08225_ _08162_ vssd1 vssd1
+ vccd1 vccd1 _08226_ sky130_fd_sc_hd__a211o_1
XFILLER_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12343_ _05525_ _05528_ _04918_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__mux2_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20413__267 clknet_1_1__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__inv_2
X_12274_ _05020_ _05458_ _05460_ _05263_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__o211a_1
X_15062_ _08156_ vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__buf_4
X_19646__28 clknet_1_1__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
XFILLER_181_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14013_ _07123_ _07122_ _07124_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__o31a_1
X_11225_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__clkinv_2
X_19870_ _03547_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11156_ _04379_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
X_18821_ _02990_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18752_ _02933_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__or2b_1
X_15964_ _09056_ _09058_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__xor2_2
X_11087_ _04343_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20559__19 clknet_1_1__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17703_ _01915_ _01990_ _01991_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__and3_1
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14915_ _08036_ _08055_ _08056_ _01633_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__o211a_1
X_18683_ _02871_ _02873_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__or2_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _08942_ _08988_ _08989_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__a21o_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _09662_ _01922_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__or3_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14846_ _07822_ _07856_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__nor2_1
X_20307__172 clknet_1_1__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__inv_2
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17565_ _10385_ _01745_ _01744_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14777_ _06655_ _07826_ _07887_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__and3_1
X_11989_ rbzero.row_render.texu\[4\] _04958_ _05042_ vssd1 vssd1 vccd1 vccd1 _05178_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_44_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19304_ rbzero.spi_registers.texadd3\[19\] _03255_ vssd1 vssd1 vccd1 vccd1 _03266_
+ sky130_fd_sc_hd__or2_1
XFILLER_72_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16516_ _09604_ _09511_ _09603_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__and3_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ _06895_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__or2b_1
XFILLER_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _08399_ _09079_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__or3_1
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19235_ rbzero.spi_registers.texadd2\[13\] _03222_ vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__or2_1
X_16447_ _09536_ _09537_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__and2b_1
XFILLER_32_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13659_ _06767_ _06808_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__nand2_1
XFILLER_176_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ rbzero.spi_registers.new_texadd\[1\]\[8\] _03174_ _03186_ _03184_ vssd1 vssd1
+ vccd1 vccd1 _00815_ sky130_fd_sc_hd__o211a_1
XFILLER_192_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16378_ _09467_ _09469_ vssd1 vssd1 vccd1 vccd1 _09470_ sky130_fd_sc_hd__nor2_1
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18117_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__or2_1
XFILLER_117_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15329_ _08144_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__nand2_1
X_19097_ rbzero.spi_registers.new_texadd\[0\]\[2\] _03141_ _03147_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00785_ sky130_fd_sc_hd__o211a_1
XFILLER_145_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03806_ _03806_ vssd1 vssd1 vccd1 vccd1 clknet_0__03806_ sky130_fd_sc_hd__clkbuf_16
X_18048_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__and2_1
XFILLER_117_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_86_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20010_ _03647_ _03650_ _03103_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__o21a_1
XFILLER_67_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19999_ _03586_ _03640_ _03641_ _03610_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__a211o_1
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21961_ net487 _01550_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ clknet_leaf_68_i_clk _00501_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21892_ net418 _01481_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ clknet_leaf_60_i_clk _00432_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20774_ rbzero.wall_tracer.rayAddendY\[-6\] _02606_ _02557_ _03956_ vssd1 vssd1 vccd1
+ vccd1 _01654_ sky130_fd_sc_hd__a22o_1
XFILLER_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_i_clk clknet_opt_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_202_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21326_ clknet_leaf_30_i_clk _00915_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21257_ clknet_leaf_0_i_clk _00846_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _04143_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20208_ rbzero.spi_registers.new_texadd\[3\]\[19\] rbzero.spi_registers.spi_buffer\[19\]
+ _03384_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
X_21188_ clknet_leaf_22_i_clk _00777_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20139_ _05650_ _09729_ _05651_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a21o_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _06124_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__nor2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _07870_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__clkbuf_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _05073_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__and2_1
X_15680_ _08246_ _08343_ _08719_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__or3_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12892_ _06058_ _06062_ _06063_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or4_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14631_ _07525_ _07579_ _07799_ _07801_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__a22oi_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _05032_ _04818_ rbzero.row_render.texu\[0\] vssd1 vssd1 vccd1 vccd1 _05033_
+ sky130_fd_sc_hd__or3b_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _10265_ _10242_ _10368_ vssd1 vssd1 vccd1 vccd1 _10369_ sky130_fd_sc_hd__a21o_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14562_ _07721_ _07732_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__xnor2_2
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _04931_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__clkbuf_8
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16301_ _08813_ _08409_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__nor2_2
XFILLER_159_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13513_ _06651_ _06609_ _06632_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__o21ai_2
X_17281_ _10160_ _10170_ _10168_ vssd1 vssd1 vccd1 vccd1 _10300_ sky130_fd_sc_hd__a21oi_1
X_10725_ _04153_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__clkbuf_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _07648_ _07662_ _07663_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__a21o_1
XFILLER_174_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19020_ _05270_ _03091_ _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__and3_4
X_16232_ _09175_ _09206_ _09324_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__a21oi_1
X_13444_ _06612_ _06614_ _06577_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__mux2_1
X_10656_ rbzero.tex_r0\[8\] rbzero.tex_r0\[7\] _04110_ vssd1 vssd1 vccd1 vccd1 _04117_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _09147_ _09149_ _09255_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__a21o_1
X_10587_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _04077_ vssd1 vssd1 vccd1 vccd1 _04081_
+ sky130_fd_sc_hd__mux2_1
X_20337__198 clknet_1_1__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__inv_2
X_13375_ _06439_ _06440_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__or2_1
XFILLER_103_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ _08207_ _08208_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__nand2_1
XFILLER_170_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ rbzero.tex_b0\[27\] _04926_ _04928_ _05198_ vssd1 vssd1 vccd1 vccd1 _05512_
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16094_ _08015_ _08018_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__or2_1
XFILLER_177_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19922_ rbzero.pov.ready_buffer\[67\] _03436_ _03582_ _08317_ _03569_ vssd1 vssd1
+ vccd1 vccd1 _03583_ sky130_fd_sc_hd__o221a_1
X_15045_ _08136_ _08140_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__nor2_1
X_12257_ rbzero.tex_g1\[41\] _04904_ _04831_ _04918_ vssd1 vssd1 vccd1 vccd1 _05444_
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11208_ _04406_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19853_ rbzero.pov.spi_buffer\[63\] rbzero.pov.spi_buffer\[64\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03539_ sky130_fd_sc_hd__mux2_1
X_12188_ _04900_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__nand2_1
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18804_ _02981_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _04370_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16996_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10017_ sky130_fd_sc_hd__or2_1
X_19784_ rbzero.pov.spi_buffer\[30\] rbzero.pov.spi_buffer\[31\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ rbzero.wall_tracer.stepDistY\[3\] _08338_ vssd1 vssd1 vccd1 vccd1 _09042_
+ sky130_fd_sc_hd__nand2_1
X_18735_ rbzero.spi_registers.spi_cmd\[2\] _02930_ rbzero.spi_registers.spi_cmd\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a21o_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18666_ _02821_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _02868_
+ sky130_fd_sc_hd__nor2_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _08930_ _08972_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__nand2_1
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17617_ _01894_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14829_ _06515_ _06498_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__nor2_2
X_18597_ rbzero.debug_overlay.vplaneY\[-5\] _02782_ vssd1 vssd1 vccd1 vccd1 _02804_
+ sky130_fd_sc_hd__or2_1
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17548_ _10094_ _01729_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__or2_1
XFILLER_205_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ _01769_ _01770_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__nor2_1
XFILLER_165_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19218_ rbzero.spi_registers.texadd2\[6\] _03208_ vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__or2_1
X_20490_ clknet_1_1__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__buf_1
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19149_ rbzero.spi_registers.new_texadd\[1\]\[0\] _03174_ _03177_ _03169_ vssd1 vssd1
+ vccd1 vccd1 _00807_ sky130_fd_sc_hd__o211a_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21111_ clknet_leaf_92_i_clk _00700_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21042_ clknet_leaf_77_i_clk _00631_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_114_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21944_ net470 _01533_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20442__293 clknet_1_1__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__inv_2
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21875_ net401 _01464_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20826_ clknet_leaf_57_i_clk _00415_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_202_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20757_ _02513_ _02518_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__and2b_1
XFILLER_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ _04038_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ rbzero.debug_overlay.playerX\[3\] vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__inv_2
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20688_ _03898_ _03901_ _03899_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__a21boi_1
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _03979_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13160_ rbzero.wall_tracer.visualWallDist\[4\] _04428_ vssd1 vssd1 vccd1 vccd1 _06331_
+ sky130_fd_sc_hd__or2_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _05299_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_21309_ clknet_leaf_35_i_clk _00898_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13091_ _06101_ _06102_ _06266_ _06265_ rbzero.wall_tracer.mapY\[6\] vssd1 vssd1
+ vccd1 vccd1 _00386_ sky130_fd_sc_hd__a32o_1
XFILLER_152_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12042_ rbzero.tex_r1\[43\] _05002_ _05230_ _04922_ vssd1 vssd1 vccd1 vccd1 _05231_
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16850_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09874_ sky130_fd_sc_hd__or2_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15801_ _08891_ _08888_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__and2b_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20525__368 clknet_1_1__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__inv_2
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16781_ _08905_ _08990_ vssd1 vssd1 vccd1 vccd1 _09813_ sky130_fd_sc_hd__and2_1
XFILLER_92_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13993_ _07150_ _07148_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__nor2_1
XFILLER_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18520_ rbzero.map_rom.f1 _02734_ _09844_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
X_15732_ _08369_ _08696_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__or2_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__clkinv_2
XFILLER_207_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _02662_ _02667_ _02677_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a21oi_1
X_15663_ _08654_ _08656_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__xnor2_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12875_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__nor2_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _10338_ _10329_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__or2b_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14614_ _07723_ _07737_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__nor2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _04958_ _05005_ _05015_ _04810_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a31o_1
X_18382_ rbzero.debug_overlay.vplaneX\[-1\] _05111_ vssd1 vssd1 vccd1 vccd1 _02614_
+ sky130_fd_sc_hd__or2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _08673_ _08686_ _08688_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__a21o_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17333_ _10328_ _10351_ vssd1 vssd1 vccd1 vccd1 _10352_ sky130_fd_sc_hd__xnor2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _07682_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__xor2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__buf_6
XFILLER_18_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ _09525_ _09243_ _10031_ _10153_ vssd1 vssd1 vccd1 vccd1 _10283_ sky130_fd_sc_hd__o31a_1
X_10708_ rbzero.tex_g1\[47\] rbzero.tex_g1\[48\] _04144_ vssd1 vssd1 vccd1 vccd1 _04145_
+ sky130_fd_sc_hd__mux2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _07592_ _07640_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__nor2_1
X_20419__273 clknet_1_0__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__inv_2
X_11688_ gpout0.hpos\[8\] _04864_ _04865_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__and3_1
XFILLER_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19003_ rbzero.spi_registers.ss_buffer\[1\] rbzero.spi_registers.ss_buffer\[0\] _03084_
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XFILLER_146_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16215_ _08012_ _08023_ _08450_ _09188_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__nor4_1
XFILLER_128_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13427_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__buf_2
X_10639_ rbzero.tex_r0\[16\] rbzero.tex_r0\[15\] _04099_ vssd1 vssd1 vccd1 vccd1 _04108_
+ sky130_fd_sc_hd__mux2_1
X_17195_ rbzero.wall_tracer.stepDistX\[8\] _09045_ _10214_ vssd1 vssd1 vccd1 vccd1
+ _10215_ sky130_fd_sc_hd__a21boi_4
XFILLER_128_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16146_ _08622_ _09082_ _09142_ _09140_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__a31o_1
X_20270__138 clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__inv_2
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _06528_ _06458_ _06459_ _06486_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__o22a_1
XFILLER_154_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ rbzero.tex_b0\[39\] _04926_ _04928_ _05198_ vssd1 vssd1 vccd1 vccd1 _05495_
+ sky130_fd_sc_hd__a31o_1
X_16077_ _09027_ _09170_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__xor2_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ _06411_ _06393_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__or2_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19905_ _08217_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__nor2_1
X_15028_ _06142_ _06248_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__nor2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19836_ rbzero.pov.spi_buffer\[55\] rbzero.pov.spi_buffer\[56\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_110_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19767_ rbzero.pov.spi_buffer\[22\] rbzero.pov.spi_buffer\[23\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16979_ _09610_ _09713_ _09712_ _09711_ vssd1 vssd1 vccd1 vccd1 _10001_ sky130_fd_sc_hd__o2bb2a_1
Xinput3 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_2
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18718_ _02914_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__nand2_1
XFILLER_188_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18649_ _02850_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__xor2_1
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21660_ clknet_leaf_17_i_clk _01249_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20611_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _03836_ vssd1 vssd1 vccd1 vccd1
+ _03841_ sky130_fd_sc_hd__a21o_1
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21591_ clknet_leaf_92_i_clk _01180_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_178_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21025_ clknet_leaf_15_i_clk _00614_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_2
XFILLER_113_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ rbzero.tex_b1\[41\] rbzero.tex_b1\[42\] _04292_ vssd1 vssd1 vccd1 vccd1 _04293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21927_ net453 _01516_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05835_ _05836_ _05838_ net23 vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__o211a_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21858_ net384 _01447_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _04748_ _04752_ _04795_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o221a_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ clknet_leaf_51_i_clk _00398_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12591_ net21 _05769_ net17 _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__and4b_1
X_21789_ net315 _01378_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _07421_ _07422_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__nand2_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _04651_ rbzero.map_overlay.i_mapdy\[1\] vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14261_ _07306_ _07203_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__or2_2
X_11473_ _04656_ rbzero.debug_overlay.playerY\[2\] vssd1 vssd1 vccd1 vccd1 _04663_
+ sky130_fd_sc_hd__or2_1
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _08628_ _08657_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__o21a_1
XFILLER_171_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13212_ rbzero.wall_tracer.visualWallDist\[-7\] _06326_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a21o_1
XFILLER_100_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10424_ _03993_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14192_ _07205_ _07210_ _07362_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__and3_1
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13143_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__or2_1
XFILLER_174_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17951_ _02237_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__and2_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _06113_ _06088_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16902_ _09921_ _09923_ vssd1 vssd1 vccd1 vccd1 _09924_ sky130_fd_sc_hd__xor2_1
X_12025_ rbzero.tex_r1\[17\] _04935_ _05186_ _04953_ vssd1 vssd1 vccd1 vccd1 _05214_
+ sky130_fd_sc_hd__a31o_1
X_17882_ _02169_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__and2_1
X_20449__299 clknet_1_1__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__inv_2
X_19621_ rbzero.pov.spi_counter\[0\] _03439_ _03441_ vssd1 vssd1 vccd1 vccd1 _01015_
+ sky130_fd_sc_hd__a21oi_1
X_16833_ _09822_ _09347_ vssd1 vssd1 vccd1 vccd1 _09859_ sky130_fd_sc_hd__nand2_1
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19552_ _03404_ vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16764_ rbzero.wall_tracer.mapX\[9\] _09119_ _09795_ vssd1 vssd1 vccd1 vccd1 _09798_
+ sky130_fd_sc_hd__o21a_1
XFILLER_20_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13976_ _07060_ _07100_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a21oi_1
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ _08710_ _08755_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__xor2_2
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18503_ rbzero.debug_overlay.playerY\[5\] _02721_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02722_ sky130_fd_sc_hd__mux2_1
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12927_ _04429_ _04430_ rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__or3b_2
XFILLER_206_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19483_ _03368_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
X_16695_ rbzero.traced_texa\[-10\] _09755_ _09754_ rbzero.wall_tracer.visualWallDist\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_94_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15646_ _08738_ _08739_ _08740_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__nand3_1
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18434_ _02597_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _02662_
+ sky130_fd_sc_hd__nand2_1
XFILLER_94_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12858_ _05995_ _06032_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__o21ai_4
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11809_ _04997_ _04998_ _04944_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__mux2_1
X_18365_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__clkbuf_4
X_15577_ _08194_ _08229_ _08233_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__or3_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12789_ _05946_ _05948_ _05962_ _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__a31o_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17316_ _10333_ _10334_ vssd1 vssd1 vccd1 vccd1 _10335_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14528_ _07693_ _07698_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__or2b_1
XFILLER_147_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18296_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__nand2_1
XFILLER_30_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _10149_ _10177_ vssd1 vssd1 vccd1 vccd1 _10266_ sky130_fd_sc_hd__nand2_1
XFILLER_186_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14459_ _07581_ _07629_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__nand2_1
X_17178_ _10196_ _10197_ vssd1 vssd1 vccd1 vccd1 _10198_ sky130_fd_sc_hd__and2b_1
XFILLER_143_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ _09089_ _09091_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__nor2_1
XFILLER_66_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ rbzero.pov.spi_buffer\[47\] rbzero.pov.spi_buffer\[48\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03521_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21712_ net238 _01301_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21643_ clknet_leaf_83_i_clk _01232_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21574_ clknet_leaf_94_i_clk _01163_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_41 _06217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22057_ clknet_leaf_40_i_clk _01646_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21008_ clknet_leaf_76_i_clk _00597_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13830_ _06992_ _06999_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__or3_1
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _06898_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__nand2_1
X_10973_ rbzero.tex_b1\[49\] rbzero.tex_b1\[50\] _04281_ vssd1 vssd1 vccd1 vccd1 _04284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15500_ _08519_ _08517_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__nand2_1
XFILLER_204_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ net33 _05887_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__and4b_1
X_16480_ _09569_ _09570_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__xnor2_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _06832_ _06833_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__nand2_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ _08496_ _08514_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__nor2_1
XFILLER_54_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ net22 vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__clkbuf_4
XFILLER_169_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18150_ _09872_ _02422_ _02337_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__o21a_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ _08456_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__buf_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12574_ _05715_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__inv_2
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17101_ _10018_ _10121_ vssd1 vssd1 vccd1 vccd1 _10122_ sky130_fd_sc_hd__xnor2_4
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14313_ _07482_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__xnor2_1
X_18081_ _02361_ _02362_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11525_ gpout0.vpos\[7\] _04713_ rbzero.map_overlay.i_otherx\[1\] _04414_ _04714_
+ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o221a_1
XFILLER_184_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15293_ _08370_ _08373_ _08386_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17032_ _10051_ _10052_ vssd1 vssd1 vccd1 vccd1 _10053_ sky130_fd_sc_hd__nor2_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14244_ _07383_ _07384_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11456_ gpout0.vpos\[3\] _04645_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__or2_1
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10407_ _03984_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14175_ _07314_ _07319_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__xor2_1
X_11387_ _04412_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__or2_1
XFILLER_113_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13126_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nor2_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ rbzero.spi_registers.spi_buffer\[22\] rbzero.spi_registers.spi_buffer\[21\]
+ _03051_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _10059_ _09621_ _02127_ _02125_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__o31a_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _06222_ _06226_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and3_1
XFILLER_26_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ rbzero.tex_r1\[7\] _05195_ _05196_ _04923_ vssd1 vssd1 vccd1 vccd1 _05197_
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20382__239 clknet_1_1__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__inv_2
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17865_ _02152_ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__nand2_1
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xnet99_2 clknet_1_0__leaf__04634_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
X_19604_ rbzero.spi_registers.new_texadd\[1\]\[19\] rbzero.spi_registers.spi_buffer\[19\]
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__mux2_1
X_16816_ _09782_ vssd1 vssd1 vccd1 vccd1 _09844_ sky130_fd_sc_hd__buf_6
X_17796_ _02085_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19535_ rbzero.spi_registers.new_texadd\[0\]\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__mux2_1
X_13959_ _07114_ _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__xnor2_2
X_16747_ _09783_ vssd1 vssd1 vccd1 vccd1 _09785_ sky130_fd_sc_hd__buf_6
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19466_ rbzero.spi_registers.new_vinf _02473_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_
+ sky130_fd_sc_hd__mux2_1
X_16678_ rbzero.row_render.size\[5\] _09746_ _09750_ _07971_ vssd1 vssd1 vccd1 vccd1
+ _00488_ sky130_fd_sc_hd__a22o_1
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18417_ _02621_ _02628_ _02629_ _02614_ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a2bb2o_1
X_15629_ _08356_ _08697_ _08699_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19397_ _02481_ rbzero.spi_registers.new_floor\[1\] _03319_ vssd1 vssd1 vccd1 vccd1
+ _03321_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18348_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__nand2_1
X_20276__144 clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__inv_2
XFILLER_159_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18279_ _02513_ _02517_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_8
XFILLER_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21290_ clknet_leaf_33_i_clk _00879_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03799_ clknet_0__03799_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03799_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20172_ _03752_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21626_ clknet_leaf_88_i_clk _01215_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21557_ clknet_leaf_90_i_clk _01146_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11310_ rbzero.texu_hot\[3\] _04484_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__or2_1
XFILLER_180_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12290_ rbzero.tex_b0\[63\] _04926_ _04928_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__and3_1
XFILLER_119_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21488_ net206 _01077_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ rbzero.trace_state\[1\] vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__buf_4
XFILLER_106_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11172_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _04384_ vssd1 vssd1 vccd1 vccd1 _04388_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15980_ _08549_ _08550_ _08552_ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__a21bo_1
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14931_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.trackDistX\[0\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__mux2_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _01718_ _01832_ _01835_ _01833_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a2bb2o_1
X_14862_ _08016_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16601_ _09690_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__buf_2
X_13813_ _06754_ _06687_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__nor2_1
XFILLER_17_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _01870_ _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__or2b_1
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14793_ _06577_ _07917_ _07903_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16532_ _08304_ _09621_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__nor2_1
X_19320_ rbzero.floor_leak\[2\] _03272_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__or2_1
XFILLER_21_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ _06913_ _06912_ _06911_ _06900_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__a211oi_1
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10956_ rbzero.tex_b1\[57\] rbzero.tex_b1\[58\] _04270_ vssd1 vssd1 vccd1 vccd1 _04275_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16463_ _09544_ _09553_ vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__xor2_2
X_19251_ rbzero.spi_registers.texadd2\[21\] _03207_ vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__or2_1
X_13675_ _06816_ _06819_ _06844_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__o211a_1
X_10887_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _04237_ vssd1 vssd1 vccd1 vccd1 _04239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _08390_ _08409_ _08384_ _08410_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__o22ai_1
X_18202_ _09872_ _02467_ _02337_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__o21a_1
X_12626_ net52 _05803_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__and2_1
X_19182_ rbzero.spi_registers.new_texadd\[1\]\[15\] _03188_ _03195_ _03184_ vssd1
+ vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__o211a_1
X_16394_ _09386_ _09403_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18133_ _02406_ _02407_ _02401_ _02403_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a211oi_1
X_15345_ _08439_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__buf_2
XFILLER_184_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12557_ _03976_ _05704_ _05703_ _05737_ net11 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a2111oi_1
XFILLER_200_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18064_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__nor2_1
X_11508_ gpout0.hpos\[2\] _04447_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__or2_1
X_15276_ _08370_ _08265_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__or2_1
XFILLER_172_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ net6 _05669_ net7 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__and3b_1
X_17015_ _09615_ _09900_ vssd1 vssd1 vccd1 vccd1 _10036_ sky130_fd_sc_hd__nand2_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14227_ _07067_ _07366_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__nand2_2
X_11439_ _04601_ _04629_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__and3_1
X_14158_ _07316_ _07303_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nor2_1
XFILLER_180_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ rbzero.wall_tracer.mapY\[10\] _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__xnor2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _03067_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__clkbuf_1
X_14089_ _06722_ _07123_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__nor2_1
XFILLER_100_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17917_ _02187_ _02204_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__xnor2_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18897_ rbzero.pov.spi_buffer\[56\] rbzero.pov.ready_buffer\[56\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
XFILLER_187_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17848_ _09670_ _01898_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__nor2_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17779_ _02066_ _02068_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__xor2_1
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19518_ rbzero.spi_registers.new_texadd\[0\]\[1\] _02481_ _03381_ vssd1 vssd1 vccd1
+ vccd1 _03387_ sky130_fd_sc_hd__mux2_1
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20790_ gpout4.clk_div\[0\] net63 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19449_ rbzero.spi_registers.got_new_other _03118_ _03316_ _03349_ vssd1 vssd1 vccd1
+ vccd1 _00935_ sky130_fd_sc_hd__a31o_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21411_ clknet_leaf_8_i_clk _01000_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21342_ clknet_leaf_9_i_clk _00931_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21273_ clknet_leaf_26_i_clk _00862_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20224_ clknet_1_0__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__buf_1
XFILLER_150_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20155_ _04731_ _03738_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nor2_1
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20086_ rbzero.debug_overlay.vplaneX\[-3\] _03685_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__or2_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _04121_ vssd1 vssd1 vccd1 vccd1 _04198_
+ sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _04978_ vssd1 vssd1 vccd1 vccd1 _04980_
+ sky130_fd_sc_hd__mux2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20988_ clknet_leaf_26_i_clk _00577_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ rbzero.tex_g1\[31\] rbzero.tex_g1\[32\] _04155_ vssd1 vssd1 vccd1 vccd1 _04162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13460_ _06537_ _06539_ _06566_ _06567_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__a31oi_4
X_10672_ _04125_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _04978_ vssd1 vssd1 vccd1 vccd1 _05596_
+ sky130_fd_sc_hd__mux2_1
X_21609_ clknet_leaf_89_i_clk _01198_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
X_13391_ _06561_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__clkinv_2
XFILLER_12_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _08220_ _06076_ _08224_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__a21oi_1
X_12342_ _05526_ _05527_ _04826_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__mux2_1
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ rbzero.trace_state\[0\] _08155_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__nand2_4
X_12273_ rbzero.row_render.texu\[2\] _04920_ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14012_ _07120_ _07121_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__nand2_1
X_11224_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__buf_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18820_ rbzero.pov.spi_buffer\[19\] rbzero.pov.ready_buffer\[19\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02990_ sky130_fd_sc_hd__mux2_1
XFILLER_96_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11155_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _04373_ vssd1 vssd1 vccd1 vccd1 _04379_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18751_ _02475_ _02932_ _02930_ rbzero.spi_registers.spi_cmd\[3\] vssd1 vssd1 vccd1
+ vccd1 _02947_ sky130_fd_sc_hd__a31o_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _08448_ _08468_ _09057_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__a21bo_1
X_11086_ rbzero.tex_b0\[60\] rbzero.tex_b0\[59\] _04340_ vssd1 vssd1 vccd1 vccd1 _04343_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17702_ _01915_ _01990_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a21oi_2
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14914_ rbzero.wall_tracer.visualWallDist\[-5\] _08047_ vssd1 vssd1 vccd1 vccd1 _08056_
+ sky130_fd_sc_hd__or2_1
X_15894_ _08906_ _08941_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__and2b_1
X_18682_ _02881_ _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nand2_1
XFILLER_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _01809_ _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14845_ _06631_ _07952_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__nand2_1
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17564_ _01771_ _01855_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__xnor2_1
X_14776_ _07903_ _07937_ _07940_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__a211oi_2
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11988_ rbzero.row_render.side _05037_ _05020_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a21o_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19303_ rbzero.spi_registers.new_texadd\[3\]\[18\] _03254_ _03264_ _03265_ vssd1
+ vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__o211a_1
XFILLER_95_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16515_ _09511_ _09603_ _09604_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__a21oi_1
X_13727_ _06895_ _06896_ _06897_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__or3_1
XFILLER_205_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10939_ rbzero.tex_g0\[2\] rbzero.tex_g0\[1\] _04259_ vssd1 vssd1 vccd1 vccd1 _04266_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17495_ _08499_ _08617_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__or2_1
XFILLER_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19234_ rbzero.spi_registers.new_texadd\[2\]\[12\] _03221_ _03225_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__o211a_1
XFILLER_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _09533_ _09535_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__nand2_1
X_13658_ _06826_ _06825_ _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__o21bai_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ net51 net41 net40 _05263_ net17 _05763_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__mux4_1
X_19165_ rbzero.spi_registers.texadd1\[8\] _03176_ vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__or2_1
X_16377_ _04686_ _09468_ _08138_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__mux2_1
XFILLER_192_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ _06681_ _06738_ _06759_ _06737_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__a22o_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15328_ _06041_ _06341_ _04464_ vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__mux2_1
X_18116_ _02393_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19096_ rbzero.spi_registers.texadd0\[2\] _03143_ vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__or2_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03805_ _03805_ vssd1 vssd1 vccd1 vccd1 clknet_0__03805_ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15259_ _08303_ _08353_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _02329_ _02333_ rbzero.wall_tracer.trackDistX\[10\] _09879_ vssd1 vssd1 vccd1
+ vccd1 _00549_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20388__245 clknet_1_0__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__inv_2
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19998_ rbzero.pov.ready_buffer\[55\] _03585_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nor2_1
XFILLER_154_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18949_ _03058_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21960_ net486 _01549_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20911_ clknet_leaf_68_i_clk _00500_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21891_ net417 _01480_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20842_ clknet_leaf_60_i_clk _00431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20773_ _02752_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21325_ clknet_leaf_29_i_clk _00914_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21256_ clknet_leaf_0_i_clk _00845_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20207_ _03770_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21187_ clknet_leaf_18_i_clk _00776_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20138_ _05651_ _05650_ _09729_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nand3_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ rbzero.pov.ready_buffer\[31\] _03687_ _03665_ vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__and3_1
X_12960_ _06125_ _06128_ _06132_ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__or4_1
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _04414_ _05075_ _05083_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__nor3_1
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\] _06065_
+ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__or4_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _07525_ _07800_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__xnor2_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11842_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14561_ _07252_ _07476_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nor2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ rbzero.tex_r0\[27\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__and3_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _09390_ _09391_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__and2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _06641_ _06576_ _06599_ _06583_ _06594_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__a32o_1
X_17280_ _10287_ _10298_ vssd1 vssd1 vccd1 vccd1 _10299_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10724_ rbzero.tex_g1\[39\] rbzero.tex_g1\[40\] _04144_ vssd1 vssd1 vccd1 vccd1 _04153_
+ sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _07649_ _07661_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__nor2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _09203_ _09205_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__and2b_1
XFILLER_110_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13443_ _06506_ _06413_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__mux2_1
X_10655_ _04116_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _09146_ _09003_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__nor2_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13374_ _06474_ _06484_ _06543_ _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__a22o_2
X_10586_ _04080_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15113_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] rbzero.debug_overlay.playerX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__o21ai_1
X_12325_ rbzero.tex_b0\[26\] _04978_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__and2_1
X_16093_ _08012_ _08015_ _08450_ _08018_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__o31a_1
XFILLER_155_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19921_ _03095_ _03436_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__nand2_1
X_15044_ _08138_ _08035_ _08139_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__a21oi_1
X_12256_ rbzero.tex_g1\[43\] _04948_ _05442_ _04827_ vssd1 vssd1 vccd1 vccd1 _05443_
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ rbzero.tex_b0\[2\] rbzero.tex_b0\[1\] _04054_ vssd1 vssd1 vccd1 vccd1 _04406_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19852_ _03538_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
X_12187_ _05019_ _05371_ _05374_ _05043_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a31o_1
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18803_ rbzero.pov.spi_buffer\[11\] rbzero.pov.ready_buffer\[11\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02981_ sky130_fd_sc_hd__mux2_1
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11138_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _04362_ vssd1 vssd1 vccd1 vccd1 _04370_
+ sky130_fd_sc_hd__mux2_1
XFILLER_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19783_ _03502_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
X_16995_ _10011_ _10016_ rbzero.wall_tracer.trackDistX\[0\] _09879_ vssd1 vssd1 vccd1
+ vccd1 _00539_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ rbzero.spi_registers.spi_cmd\[0\] rbzero.spi_registers.spi_cmd\[1\] vssd1
+ vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__or2_2
X_15946_ _09039_ _09040_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__xnor2_2
X_11069_ rbzero.tex_b1\[3\] rbzero.tex_b1\[4\] _04325_ vssd1 vssd1 vccd1 vccd1 _04334_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ _02847_ _02853_ _02841_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a21o_1
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _08928_ _08929_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__or2_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20502__347 clknet_1_0__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__inv_2
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17616_ _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__nor2_1
X_14828_ _07826_ _07986_ _07987_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__a21bo_1
X_18596_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nand2_1
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ _10221_ _01729_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__nand2_1
X_14759_ _07854_ _07925_ _07827_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__mux2_1
XFILLER_177_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17478_ _01689_ _01767_ _01768_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__and3_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19217_ rbzero.spi_registers.new_texadd\[2\]\[5\] _03206_ _03216_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00836_ sky130_fd_sc_hd__o211a_1
X_16429_ _08734_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19148_ rbzero.spi_registers.texadd1\[0\] _03176_ vssd1 vssd1 vccd1 vccd1 _03177_
+ sky130_fd_sc_hd__or2_1
XFILLER_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19079_ rbzero.mapdxw\[0\] _03121_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or2_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21110_ clknet_leaf_92_i_clk _00699_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21041_ clknet_leaf_86_i_clk _00630_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21943_ net469 _01532_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21874_ net400 _01463_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ clknet_leaf_58_i_clk _00414_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20756_ rbzero.wall_tracer.rayAddendX\[-8\] _02606_ _02557_ _03944_ vssd1 vssd1 vccd1
+ vccd1 _01648_ sky130_fd_sc_hd__a22o_1
XFILLER_195_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20687_ _03903_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__and2b_1
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _04001_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ reg_rgb\[7\] _05298_ _05058_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__mux2_4
X_21308_ clknet_leaf_35_i_clk _00897_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ _06105_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__nor2_2
XFILLER_123_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12041_ rbzero.tex_r1\[42\] _05031_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__or2_1
X_21239_ clknet_leaf_4_i_clk _00828_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _08870_ _08894_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__or2_1
XFILLER_120_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16780_ _09782_ vssd1 vssd1 vccd1 vccd1 _09812_ sky130_fd_sc_hd__buf_4
XFILLER_19_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13992_ _07145_ _07147_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__nor2_1
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15731_ _08821_ _08825_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__xor2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ rbzero.debug_overlay.playerX\[1\] _06117_ _06080_ rbzero.debug_overlay.playerY\[5\]
+ _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a221o_1
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _02597_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 _02677_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15662_ _08756_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__inv_2
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _06010_ _06017_ _06005_ rbzero.wall_tracer.rayAddendY\[3\] rbzero.debug_overlay.facingY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a32o_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _10317_ _10325_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_85_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _04941_ _05008_ _05014_ _04955_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a211o_1
X_14613_ _07780_ _07768_ _07781_ _07782_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_2_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15593_ _08687_ _08299_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__xor2_1
X_18381_ _02610_ _02611_ _02608_ _02609_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a211o_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17332_ _10348_ _10350_ vssd1 vssd1 vccd1 vccd1 _10351_ sky130_fd_sc_hd__xnor2_1
X_14544_ _07708_ _07707_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__and2b_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _04826_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__buf_4
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17263_ _10280_ _10281_ vssd1 vssd1 vccd1 vccd1 _10282_ sky130_fd_sc_hd__or2_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _07603_ _07616_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11687_ _03972_ _04867_ _04868_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a22o_1
XFILLER_201_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19002_ _03086_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16214_ _09053_ _09306_ _08441_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__a21oi_2
X_13426_ _06569_ _06538_ _06570_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__and3_1
X_10638_ _04107_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__clkbuf_1
X_17194_ _06263_ _09426_ vssd1 vssd1 vccd1 vccd1 _10214_ sky130_fd_sc_hd__nand2_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _09227_ _09228_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__nand2_1
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13357_ _06344_ _06450_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__xnor2_1
X_10569_ _04071_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ rbzero.tex_b0\[38\] _05314_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__and2_1
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ _08369_ _08497_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_23_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13288_ _06451_ _06455_ _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__or3_2
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19904_ _03437_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__buf_2
XFILLER_64_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15027_ _08124_ _08033_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__nand2_1
XFILLER_170_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ rbzero.tex_g1\[49\] _04904_ _04831_ _04918_ vssd1 vssd1 vccd1 vccd1 _05426_
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19835_ _03529_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19766_ _03493_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16978_ _09998_ _09999_ vssd1 vssd1 vccd1 vccd1 _10000_ sky130_fd_sc_hd__nand2_1
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
X_18717_ _02822_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _02915_
+ sky130_fd_sc_hd__nand2_1
X_15929_ _09001_ _09023_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18648_ _02833_ _02838_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__or2b_1
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18579_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__nand2_1
XFILLER_33_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20610_ _03838_ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2b_1
XFILLER_178_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21590_ clknet_leaf_15_i_clk _01179_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__05938_ _05938_ vssd1 vssd1 vccd1 vccd1 clknet_0__05938_ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22073_ clknet_leaf_38_i_clk _01662_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21024_ clknet_leaf_15_i_clk _00613_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_2
XFILLER_102_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21926_ net452 _01515_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21857_ net383 _01446_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11610_ _04751_ _04796_ _04797_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o21ai_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20808_ clknet_leaf_51_i_clk _00397_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12590_ net18 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__buf_2
X_21788_ net314 _01377_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _04656_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__inv_2
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20739_ rbzero.traced_texVinit\[4\] _09759_ _03937_ _09347_ vssd1 vssd1 vccd1 vccd1
+ _01638_ sky130_fd_sc_hd__a22o_1
XFILLER_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _07429_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__nand2_1
XFILLER_184_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _04656_ rbzero.debug_overlay.playerY\[2\] vssd1 vssd1 vccd1 vccd1 _04662_
+ sky130_fd_sc_hd__nand2_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13211_ _06380_ _06381_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__xor2_4
X_10423_ rbzero.tex_r1\[52\] rbzero.tex_r1\[53\] _03991_ vssd1 vssd1 vccd1 vccd1 _03993_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14191_ _06720_ _07361_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__nor2_1
XFILLER_139_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__nand2_1
XFILLER_87_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17950_ _02235_ _02236_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__nand2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _06144_ rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16901_ _09626_ _09631_ _09922_ vssd1 vssd1 vccd1 vccd1 _09923_ sky130_fd_sc_hd__a21boi_1
X_12024_ rbzero.tex_r1\[19\] _04933_ _05212_ _05191_ vssd1 vssd1 vccd1 vccd1 _05213_
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17881_ _02167_ _02168_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__nand2_1
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19620_ rbzero.pov.spi_counter\[0\] _03439_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_
+ sky130_fd_sc_hd__o21ai_1
X_16832_ _09854_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09858_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19551_ rbzero.spi_registers.new_texadd\[0\]\[17\] rbzero.spi_registers.spi_buffer\[17\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16763_ rbzero.wall_tracer.mapX\[9\] _09786_ _09784_ _09797_ vssd1 vssd1 vccd1 vccd1
+ _00526_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13975_ _07063_ _07099_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__and2b_1
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18502_ _06081_ _02720_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _08765_ _08808_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__nor2_1
XFILLER_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12926_ _06100_ _06079_ _06099_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or3_1
X_19482_ rbzero.spi_registers.new_mapd\[5\] _02489_ _03362_ vssd1 vssd1 vccd1 vccd1
+ _03368_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16694_ _09751_ vssd1 vssd1 vccd1 vccd1 _09755_ sky130_fd_sc_hd__clkbuf_4
XFILLER_62_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18433_ _02661_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15645_ _08668_ _08730_ _08737_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__a21o_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12857_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__or2_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _04909_ vssd1 vssd1 vccd1 vccd1 _04998_
+ sky130_fd_sc_hd__mux2_1
X_18364_ _02596_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__buf_2
X_15576_ _08227_ _08252_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__or2_1
X_12788_ _05963_ _05964_ _05948_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__mux2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17315_ _08889_ _09680_ vssd1 vssd1 vccd1 vccd1 _10334_ sky130_fd_sc_hd__and2b_1
X_11739_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__buf_4
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14527_ _07693_ _07695_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__or3_2
X_18295_ _08135_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17246_ _10239_ _10240_ vssd1 vssd1 vccd1 vccd1 _10265_ sky130_fd_sc_hd__or2_1
X_14458_ _06857_ _07209_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _06577_ _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__xnor2_4
X_17177_ _10193_ _10195_ vssd1 vssd1 vccd1 vccd1 _10197_ sky130_fd_sc_hd__nand2_1
X_14389_ _07508_ _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__nand2_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16128_ _09086_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__xnor2_4
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16059_ _09151_ _09152_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20508__353 clknet_1_1__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__inv_2
X_19818_ _03520_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19749_ _03484_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21711_ net237 _01300_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21642_ clknet_leaf_83_i_clk _01231_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_20 rbzero.tex_r0\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21573_ clknet_leaf_94_i_clk _01162_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_42 _07996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20253__123 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__inv_2
XFILLER_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19693__71 clknet_1_0__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_121_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22056_ clknet_leaf_40_i_clk _01645_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21007_ clknet_leaf_79_i_clk _00596_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _06895_ _06896_ _06897_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__o21ai_1
X_10972_ _04283_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21909_ net435 _01498_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
X_12711_ net30 vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__buf_2
XFILLER_189_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13691_ _06853_ _06861_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__xnor2_2
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12642_ _05821_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
X_15430_ _08520_ _08524_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ rbzero.wall_tracer.visualWallDist\[-10\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _08456_ sky130_fd_sc_hd__nand2_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ net53 _05720_ _05715_ net55 _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a221o_1
XFILLER_196_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ _09894_ _10120_ vssd1 vssd1 vccd1 vccd1 _10121_ sky130_fd_sc_hd__xnor2_4
XFILLER_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14312_ _07115_ _07309_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__and2_1
X_11524_ _04648_ rbzero.map_overlay.i_othery\[3\] vssd1 vssd1 vccd1 vccd1 _04714_
+ sky130_fd_sc_hd__xnor2_1
X_15292_ _08370_ _08373_ _08386_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__or3_1
X_18080_ _02353_ _02355_ _02354_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a21boi_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17031_ _10049_ _10050_ vssd1 vssd1 vccd1 vccd1 _10052_ sky130_fd_sc_hd__and2_1
X_14243_ _07380_ _07388_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__xnor2_1
X_11455_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__or2_1
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ rbzero.tex_r1\[60\] rbzero.tex_r1\[61\] _03980_ vssd1 vssd1 vccd1 vccd1 _03984_
+ sky130_fd_sc_hd__mux2_1
X_14174_ _07115_ _07331_ _07344_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a21o_1
XFILLER_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13125_ _06292_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nand2_1
XFILLER_113_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18982_ _03075_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _02219_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nand2_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _06223_ _06227_ _06230_ _06231_ _06158_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__o2111a_1
XFILLER_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ rbzero.tex_r1\[6\] _05182_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__or2_1
X_17864_ _02122_ _02123_ _02151_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__nand3_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19603_ _03430_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__clkbuf_1
X_16815_ _09839_ _09840_ _09841_ _06104_ vssd1 vssd1 vccd1 vccd1 _09843_ sky130_fd_sc_hd__a31o_1
XFILLER_113_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ rbzero.wall_tracer.trackDistX\[7\] _02084_ _09844_ vssd1 vssd1 vccd1 vccd1
+ _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19534_ _03380_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__buf_4
X_16746_ _06105_ _09783_ vssd1 vssd1 vccd1 vccd1 _09784_ sky130_fd_sc_hd__nor2_2
X_13958_ _07127_ _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__and2_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19465_ _02474_ _08116_ _03350_ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1
+ vccd1 _03358_ sky130_fd_sc_hd__and4b_1
X_12909_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__inv_2
X_16677_ rbzero.row_render.size\[4\] _09746_ _09750_ _07964_ vssd1 vssd1 vccd1 vccd1
+ _00487_ sky130_fd_sc_hd__a22o_1
XFILLER_185_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13889_ _06779_ _06884_ _07059_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__a21bo_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18416_ _02644_ _02645_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__nor2_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ _08717_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__or2b_1
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19396_ _03320_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18347_ _02581_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15559_ _08629_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__xor2_1
XFILLER_187_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18278_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__nand2_1
X_17229_ _10006_ _10122_ vssd1 vssd1 vccd1 vccd1 _10249_ sky130_fd_sc_hd__nand2_1
Xinput40 i_mode[0] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_16
XFILLER_147_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput51 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_8
XFILLER_175_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03798_ clknet_0__03798_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03798_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20171_ rbzero.spi_registers.new_texadd\[3\]\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__mux2_1
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21625_ clknet_leaf_87_i_clk _01214_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21556_ clknet_leaf_13_i_clk _01145_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21487_ net205 _01076_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11240_ rbzero.trace_state\[3\] _04429_ _04430_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_
+ sky130_fd_sc_hd__o31a_1
XFILLER_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ _04387_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22039_ clknet_leaf_34_i_clk _01628_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14930_ _08065_ _08066_ _08067_ _08061_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__o211a_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ rbzero.wall_tracer.stepDistY\[5\] _08015_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08016_ sky130_fd_sc_hd__mux2_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16600_ _08039_ _08338_ _09689_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__or3_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _06982_ _06726_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__or2_1
XFILLER_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17580_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__nand2_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14792_ _07894_ _07909_ _07912_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__a21o_1
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16531_ _09491_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__buf_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10955_ _04274_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
X_13743_ _06900_ _06911_ _06912_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__o211a_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19250_ rbzero.spi_registers.new_texadd\[2\]\[20\] _03205_ _03234_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__o211a_1
XFILLER_189_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16462_ _09546_ _09552_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__xor2_2
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ _04238_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
X_13674_ _06827_ _06843_ _06829_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__nand3_1
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ _02464_ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__xnor2_1
X_15413_ _08410_ _08408_ _08507_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__or3b_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ net46 _05802_ _05803_ net43 _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a221o_1
X_19181_ rbzero.spi_registers.texadd1\[15\] _03189_ vssd1 vssd1 vccd1 vccd1 _03195_
+ sky130_fd_sc_hd__or2_1
X_16393_ _09379_ _09380_ _09381_ _09367_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18132_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nand2_1
XFILLER_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15344_ rbzero.wall_tracer.visualWallDist\[-9\] _06260_ _08162_ rbzero.debug_overlay.playerX\[-9\]
+ _08438_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__a221oi_2
X_12556_ _03975_ _05704_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nor2_1
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ gpout0.vpos\[9\] _04420_ net1 vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__or3b_1
XFILLER_172_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18063_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ _02344_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15275_ _08201_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__clkbuf_4
X_12487_ net41 _05664_ _05663_ _05263_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a221o_1
XFILLER_144_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ _10033_ _10034_ vssd1 vssd1 vccd1 vccd1 _10035_ sky130_fd_sc_hd__xnor2_1
X_14226_ _07331_ _07396_ _07333_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__or3b_1
X_11438_ _04410_ _04423_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__xnor2_2
X_14157_ _07306_ _07305_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__or2_1
X_11369_ rbzero.spi_registers.texadd3\[22\] _04526_ _04560_ vssd1 vssd1 vccd1 vccd1
+ _04561_ sky130_fd_sc_hd__a21o_1
XFILLER_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13108_ rbzero.wall_tracer.mapY\[9\] _06078_ _06279_ vssd1 vssd1 vccd1 vccd1 _06280_
+ sky130_fd_sc_hd__a21oi_1
X_19672__52 clknet_1_1__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ rbzero.spi_registers.spi_buffer\[13\] rbzero.spi_registers.spi_buffer\[12\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
X_14088_ _07178_ _07222_ _07233_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _02202_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nor2_1
XFILLER_117_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _06164_ rbzero.wall_tracer.trackDistY\[10\] _06214_ vssd1 vssd1 vccd1 vccd1
+ _06215_ sky130_fd_sc_hd__o21a_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ _03029_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17847_ _01923_ _02044_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__nand2_1
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17778_ _01918_ _01957_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19517_ _03386_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__clkbuf_1
X_16729_ rbzero.map_rom.f4 _09766_ vssd1 vssd1 vccd1 vccd1 _09767_ sky130_fd_sc_hd__and2_1
XFILLER_207_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19448_ _03338_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__inv_2
XFILLER_210_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19379_ _03310_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20471__319 clknet_1_0__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__inv_2
XFILLER_124_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21410_ clknet_leaf_7_i_clk _00999_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21341_ clknet_leaf_8_i_clk _00930_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21272_ clknet_leaf_25_i_clk _00861_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20154_ _04731_ _03738_ _03739_ _03740_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a211oi_1
X_20365__224 clknet_1_1__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__inv_2
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20085_ rbzero.debug_overlay.vplaneX\[-4\] _03676_ _03696_ _03695_ vssd1 vssd1 vccd1
+ vccd1 _01224_ sky130_fd_sc_hd__a211o_1
XFILLER_44_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20987_ clknet_leaf_26_i_clk _00576_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ _04161_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _04121_ vssd1 vssd1 vccd1 vccd1 _04125_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _05593_ _05594_ _05190_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__mux2_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21608_ clknet_leaf_88_i_clk _01197_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13390_ _06474_ _06508_ _06510_ _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__or4_1
XFILLER_90_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _04892_ vssd1 vssd1 vccd1 vccd1 _05527_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21539_ clknet_leaf_73_i_clk _01128_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ rbzero.trace_state\[1\] _06259_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__and2_1
XFILLER_181_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ rbzero.row_render.texu\[2\] _04920_ _05019_ vssd1 vssd1 vccd1 vccd1 _05459_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ _07089_ _07090_ _07137_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__and3_1
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__clkbuf_4
XFILLER_181_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _04378_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18750_ rbzero.spi_registers.spi_counter\[4\] _02934_ _02945_ vssd1 vssd1 vccd1 vccd1
+ _02946_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15962_ _09043_ _08581_ _08467_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__or3_1
X_11085_ _04342_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17701_ _01891_ _01892_ _01889_ _01890_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14913_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.trackDistX\[-5\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__mux2_1
X_18681_ rbzero.debug_overlay.vplaneY\[-2\] _02868_ vssd1 vssd1 vccd1 vccd1 _02882_
+ sky130_fd_sc_hd__nand2_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _08868_ _08983_ _08985_ _08987_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__and4_1
XFILLER_23_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _01697_ _09315_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__nor2_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ _08001_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17563_ _01852_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__xor2_1
XFILLER_189_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _06633_ _06602_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__nand2_1
XFILLER_44_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11987_ _04589_ _05061_ _05063_ _05175_ _04650_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__o311a_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19302_ _03212_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__buf_4
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _09487_ _09494_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__or2b_1
XFILLER_32_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _06726_ _06798_ _06700_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
X_10938_ _04265_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17494_ _01702_ _01703_ _01698_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__o21ai_1
XFILLER_210_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19709__86 clknet_1_1__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19233_ _03212_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__clkbuf_4
X_16445_ _09533_ _09535_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__nor2_1
X_10869_ _04229_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
X_13657_ _06736_ _06740_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__nand2_1
XFILLER_32_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _05772_ _05787_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__and4b_1
X_19164_ rbzero.spi_registers.new_texadd\[1\]\[7\] _03174_ _03185_ _03184_ vssd1 vssd1
+ vccd1 vccd1 _00814_ sky130_fd_sc_hd__o211a_1
XFILLER_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__clkinv_2
X_13588_ _06708_ _06734_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and2_2
XFILLER_30_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18115_ rbzero.wall_tracer.trackDistY\[-3\] _02392_ _02339_ vssd1 vssd1 vccd1 vccd1
+ _02393_ sky130_fd_sc_hd__mux2_1
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15327_ rbzero.wall_tracer.stepDistY\[1\] vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__inv_2
X_19095_ rbzero.spi_registers.new_texadd\[0\]\[1\] _03141_ _03146_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00784_ sky130_fd_sc_hd__o211a_1
X_12539_ _05702_ _05704_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__and2_1
XFILLER_144_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03804_ _03804_ vssd1 vssd1 vccd1 vccd1 clknet_0__03804_ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18046_ _08124_ _02332_ _09783_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a21oi_1
X_15258_ _08306_ _08352_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14209_ _07363_ _07379_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__xor2_1
X_20314__178 clknet_1_0__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__inv_2
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15189_ _08283_ rbzero.debug_overlay.playerY\[-3\] _06076_ vssd1 vssd1 vccd1 vccd1
+ _08284_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19997_ rbzero.debug_overlay.playerY\[2\] rbzero.debug_overlay.playerY\[1\] _03632_
+ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__or3_1
XFILLER_67_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18948_ _02489_ _02487_ _03052_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
XFILLER_79_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18879_ _03020_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20910_ clknet_leaf_50_i_clk _00499_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
X_21890_ net416 _01479_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20841_ clknet_leaf_60_i_clk _00430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20772_ _05129_ rbzero.wall_tracer.rayAddendY\[-6\] vssd1 vssd1 vccd1 vccd1 _03955_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21324_ clknet_leaf_30_i_clk _00913_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21255_ clknet_leaf_1_i_clk _00844_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20206_ rbzero.spi_registers.new_texadd\[3\]\[18\] rbzero.spi_registers.spi_buffer\[18\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__mux2_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21186_ clknet_leaf_18_i_clk _00775_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20137_ _08116_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__clkbuf_4
X_19651__33 clknet_1_0__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _03096_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__buf_2
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20549__10 clknet_1_1__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _05095_ _05096_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__or3_1
XFILLER_206_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__xor2_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _04829_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__clkbuf_4
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20564__24 clknet_1_0__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11772_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _04914_ vssd1 vssd1 vccd1 vccd1 _04962_
+ sky130_fd_sc_hd__mux2_1
X_14560_ _07696_ _07727_ _07728_ _07730_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__a22o_2
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _04152_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__clkbuf_1
X_13511_ _06658_ _06671_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a21o_4
XFILLER_53_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14491_ _07649_ _07661_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__xor2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16230_ _09301_ _09322_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__xnor2_1
X_10654_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _04110_ vssd1 vssd1 vccd1 vccd1 _04116_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13442_ _06590_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16161_ _09251_ _09253_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__nand2_1
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13373_ _06480_ _06514_ _06448_ _06467_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__and4bb_2
X_10585_ rbzero.tex_r0\[42\] rbzero.tex_r0\[41\] _04077_ vssd1 vssd1 vccd1 vccd1 _04080_
+ sky130_fd_sc_hd__mux2_1
XFILLER_177_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15112_ rbzero.debug_overlay.playerX\[-7\] rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__or3_1
X_12324_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _04908_ vssd1 vssd1 vccd1 vccd1 _05510_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16092_ _09185_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__buf_2
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12255_ rbzero.tex_g1\[42\] _04829_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__or2_1
X_19920_ rbzero.debug_overlay.playerX\[-2\] _03569_ _03581_ _03579_ vssd1 vssd1 vccd1
+ vccd1 _01174_ sky130_fd_sc_hd__o211a_1
X_15043_ _06217_ _08035_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__nor2_1
XFILLER_135_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11206_ _04405_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19851_ rbzero.pov.spi_buffer\[62\] rbzero.pov.spi_buffer\[63\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_1
X_12186_ rbzero.row_render.side _05033_ _05373_ _05038_ _05020_ vssd1 vssd1 vccd1
+ vccd1 _05374_ sky130_fd_sc_hd__a311o_1
XFILLER_123_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11137_ _04369_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18802_ _02980_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19782_ rbzero.pov.spi_buffer\[29\] rbzero.pov.spi_buffer\[30\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XFILLER_150_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16994_ _09872_ _10014_ _10015_ _09879_ vssd1 vssd1 vccd1 vccd1 _10016_ sky130_fd_sc_hd__o31a_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__buf_2
X_15945_ _08434_ _08497_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__nor2_1
X_11068_ _04333_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18664_ _02863_ _02864_ _02862_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21o_1
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _08949_ _08956_ _08959_ _08969_ _08970_ vssd1 vssd1 vccd1 vccd1 _08971_ sky130_fd_sc_hd__a311o_1
XFILLER_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17615_ _01895_ _01896_ _01904_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__and3_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14827_ _06595_ _07959_ _07960_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__or3_1
X_18595_ _02800_ _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__nand2_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17546_ _01830_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__xnor2_1
X_14758_ _07848_ _07857_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13709_ _06770_ _06877_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__or2_1
X_17477_ _01689_ _01767_ _01768_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a21oi_1
XFILLER_204_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14689_ _06613_ _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__nor2_1
X_20394__250 clknet_1_1__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__inv_2
XFILLER_60_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19216_ rbzero.spi_registers.texadd2\[5\] _03208_ vssd1 vssd1 vccd1 vccd1 _03216_
+ sky130_fd_sc_hd__or2_1
X_16428_ _08666_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19147_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__buf_2
X_16359_ _09449_ _09450_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__and2b_1
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19078_ rbzero.spi_registers.new_mapd\[9\] _03119_ _03135_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00778_ sky130_fd_sc_hd__o211a_1
XFILLER_69_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18029_ _02314_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21040_ clknet_leaf_78_i_clk _00629_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_158_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21942_ net468 _01531_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21873_ net399 _01462_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20477__325 clknet_1_1__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__inv_2
X_20824_ clknet_leaf_58_i_clk _00413_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20755_ _02514_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20686_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _03904_
+ sky130_fd_sc_hd__nand2_1
XFILLER_206_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21307_ clknet_leaf_30_i_clk _00896_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12040_ rbzero.tex_r1\[44\] _04935_ _05195_ _05227_ _05228_ vssd1 vssd1 vccd1 vccd1
+ _05229_ sky130_fd_sc_hd__a311o_1
XFILLER_3_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21238_ clknet_leaf_4_i_clk _00827_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21169_ clknet_leaf_9_i_clk _00758_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13991_ _07148_ _07151_ _07153_ _07108_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15730_ _08822_ _08824_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__xnor2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _06111_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__nor2_1
XFILLER_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _08710_ _08755_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__nor2_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12873_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__or2_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17400_ _10322_ _10324_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__nor2_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07780_ _07768_ _07781_ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11824_ _05011_ _05012_ _05013_ _04947_ _04919_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__o221a_1
X_18380_ _02608_ _02609_ _02610_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__o211ai_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08300_ _08291_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__nand2_1
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _10213_ _10223_ _10349_ vssd1 vssd1 vccd1 vccd1 _10350_ sky130_fd_sc_hd__a21bo_1
XFILLER_144_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07674_ _07712_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__xor2_1
X_11755_ _04942_ _04943_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__mux2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _10278_ _10279_ vssd1 vssd1 vccd1 vccd1 _10281_ sky130_fd_sc_hd__nor2_1
X_10706_ _03978_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__buf_4
XFILLER_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14474_ _07642_ _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__nor2_1
X_11686_ _04874_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand2_1
XFILLER_202_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19001_ net43 rbzero.spi_registers.ss_buffer\[0\] _09734_ vssd1 vssd1 vccd1 vccd1
+ _03086_ sky130_fd_sc_hd__mux2_1
X_16213_ rbzero.wall_tracer.stepDistX\[5\] _09045_ vssd1 vssd1 vccd1 vccd1 _09306_
+ sky130_fd_sc_hd__nand2_4
X_13425_ _06583_ _06593_ _06595_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__mux2_1
X_10637_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _04099_ vssd1 vssd1 vccd1 vccd1 _04107_
+ sky130_fd_sc_hd__mux2_1
X_17193_ _10203_ _10212_ vssd1 vssd1 vccd1 vccd1 _10213_ sky130_fd_sc_hd__xor2_1
XFILLER_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ rbzero.texu_hot\[1\] _08145_ _09237_ _08085_ vssd1 vssd1 vccd1 vccd1 _00467_
+ sky130_fd_sc_hd__o211a_1
X_10568_ rbzero.tex_r0\[50\] rbzero.tex_r0\[49\] _04066_ vssd1 vssd1 vccd1 vccd1 _04071_
+ sky130_fd_sc_hd__mux2_1
X_13356_ _06516_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__or2_1
XFILLER_143_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _04908_ vssd1 vssd1 vccd1 vccd1 _05493_
+ sky130_fd_sc_hd__mux2_1
X_16075_ _09167_ _08497_ _09039_ _09168_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__o31a_1
XFILLER_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10499_ _04032_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13287_ _06456_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__xor2_2
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15026_ _08123_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__buf_6
XFILLER_29_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19903_ _03565_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__clkbuf_4
X_12238_ rbzero.tex_g1\[51\] _04948_ _05424_ _04827_ vssd1 vssd1 vccd1 vccd1 _05425_
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12169_ rbzero.tex_g0\[51\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__and3_1
X_19834_ rbzero.pov.spi_buffer\[54\] rbzero.pov.spi_buffer\[55\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03529_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16977_ _09896_ _09997_ vssd1 vssd1 vccd1 vccd1 _09999_ sky130_fd_sc_hd__or2_1
X_19765_ rbzero.pov.spi_buffer\[21\] rbzero.pov.spi_buffer\[22\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03493_ sky130_fd_sc_hd__mux2_1
XFILLER_84_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_6
XFILLER_209_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ _09021_ _09022_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__nand2_1
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18716_ _02822_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__or2_1
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20426__279 clknet_1_0__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__inv_2
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18647_ _05127_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _02850_
+ sky130_fd_sc_hd__xor2_1
X_15859_ _08296_ _08473_ _08458_ _08335_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__o22a_1
XFILLER_25_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18578_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__or2_1
XFILLER_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ _10318_ _01705_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__nand2_1
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22072_ clknet_leaf_38_i_clk _01661_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21023_ clknet_leaf_15_i_clk _00612_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_1
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21925_ net451 _01514_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21856_ net382 _01445_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20807_ clknet_leaf_51_i_clk _00396_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21787_ net313 _01376_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11540_ rbzero.map_overlay.i_mapdy\[3\] vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__inv_2
X_20738_ rbzero.traced_texVinit\[3\] _09759_ _03937_ _09227_ vssd1 vssd1 vccd1 vccd1
+ _01637_ sky130_fd_sc_hd__a22o_1
XFILLER_195_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11471_ _04650_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and2_1
X_20669_ _03883_ _03886_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nand2_1
XFILLER_11_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _03992_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__clkbuf_1
X_13210_ _06298_ _06301_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__and2b_1
XFILLER_100_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_178_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20531__374 clknet_1_0__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__inv_2
XFILLER_3_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13141_ _06311_ _06290_ _06289_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20230__102 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__inv_2
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13072_ _04705_ rbzero.map_rom.f2 _06236_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16900_ _09625_ _09632_ vssd1 vssd1 vccd1 vccd1 _09922_ sky130_fd_sc_hd__nand2_1
X_12023_ rbzero.tex_r1\[18\] _05182_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__or2_1
XFILLER_151_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17880_ _02167_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__or2_1
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16831_ _09854_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09857_ sky130_fd_sc_hd__and3_1
XFILLER_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19550_ _03403_ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16762_ _09795_ _09796_ vssd1 vssd1 vccd1 vccd1 _09797_ sky130_fd_sc_hd__xnor2_1
X_13974_ _07110_ _07144_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__xor2_1
XFILLER_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18501_ rbzero.map_rom.i_row\[4\] _06078_ _06098_ vssd1 vssd1 vccd1 vccd1 _02720_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_185_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15713_ _08782_ _08806_ _08807_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19481_ _03367_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
X_12925_ _06079_ _06099_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16693_ rbzero.traced_texa\[-11\] _09752_ _09754_ rbzero.wall_tracer.visualWallDist\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
XFILLER_206_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18432_ rbzero.wall_tracer.rayAddendX\[6\] _02660_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02661_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15644_ _08714_ _08713_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__xor2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05996_ _05998_ _06029_ _06030_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a41o_2
XFILLER_181_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _04909_ vssd1 vssd1 vccd1 vccd1 _04997_
+ sky130_fd_sc_hd__mux2_1
X_18363_ rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__buf_2
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _08639_ _08664_ _08669_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__nand3_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _04420_ _05944_ _05941_ _03975_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a22o_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17314_ _08816_ _09559_ vssd1 vssd1 vccd1 vccd1 _10333_ sky130_fd_sc_hd__nor2_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _06959_ _07248_ _07696_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__o21ba_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11738_ _04828_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__clkbuf_4
X_18294_ _02531_ _02532_ _08136_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ _10135_ _10139_ _10261_ _10262_ vssd1 vssd1 vccd1 vccd1 _10264_ sky130_fd_sc_hd__a211oi_2
X_14457_ _07598_ _07622_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__xnor2_1
X_19679__58 clknet_1_1__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
X_11669_ _04412_ _04852_ _04850_ gpout0.hpos\[4\] _04858_ vssd1 vssd1 vccd1 vccd1
+ _04859_ sky130_fd_sc_hd__a221o_1
XFILLER_190_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13408_ _06578_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__buf_4
X_17176_ _10193_ _10195_ vssd1 vssd1 vccd1 vccd1 _10196_ sky130_fd_sc_hd__nor2_1
XFILLER_190_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14388_ _06757_ _07417_ _07303_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ _09219_ _09220_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__and2b_1
XFILLER_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13339_ _06391_ _06509_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__xnor2_4
XFILLER_116_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16058_ _08368_ _08328_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__nor2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ _08114_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19817_ rbzero.pov.spi_buffer\[46\] rbzero.pov.spi_buffer\[47\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03520_ sky130_fd_sc_hd__mux2_1
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19748_ rbzero.pov.spi_buffer\[13\] rbzero.pov.spi_buffer\[14\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_38_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21710_ net236 _01299_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ clknet_leaf_80_i_clk _01230_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21572_ clknet_leaf_94_i_clk _01161_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
XANTENNA_10 _08039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20523_ clknet_1_0__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__buf_1
XFILLER_162_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_43 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_84_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22055_ clknet_leaf_54_i_clk _01644_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21006_ clknet_leaf_25_i_clk _00595_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_99_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_210_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10971_ rbzero.tex_b1\[50\] rbzero.tex_b1\[51\] _04281_ vssd1 vssd1 vccd1 vccd1 _04283_
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ net29 vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__buf_2
X_21908_ net434 _01497_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13690_ _06855_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xnor2_2
XFILLER_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12641_ reg_gpout\[2\] clknet_1_1__leaf__05820_ net45 vssd1 vssd1 vccd1 vccd1 _05821_
+ sky130_fd_sc_hd__mux2_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21839_ net365 _01428_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15360_ _08148_ _08450_ _08451_ _08454_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__a31o_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ net52 _05719_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__and2_1
XFILLER_184_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _07045_ _07366_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__nor2_1
X_11523_ rbzero.map_overlay.i_othery\[4\] vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__inv_2
XFILLER_184_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15291_ _08377_ _08385_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_37_i_clk clknet_opt_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ _10049_ _10050_ vssd1 vssd1 vccd1 vccd1 _10051_ sky130_fd_sc_hd__nor2_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _07392_ _07391_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__xor2_2
X_11454_ gpout0.vpos\[9\] gpout0.vpos\[8\] _04642_ _04643_ vssd1 vssd1 vccd1 vccd1
+ _04644_ sky130_fd_sc_hd__or4_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _03983_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14173_ _07252_ _07303_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__nor2_1
X_11385_ _04449_ _04571_ _04572_ _04576_ _04446_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a311o_1
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ _06293_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__or2b_1
X_18981_ rbzero.spi_registers.spi_buffer\[21\] rbzero.spi_registers.spi_buffer\[20\]
+ _03051_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XFILLER_113_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17932_ _10315_ _09621_ _02218_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__o21ai_1
XFILLER_139_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ rbzero.map_rom.f4 rbzero.map_rom.f2 _06088_ rbzero.map_rom.b6 vssd1 vssd1
+ vccd1 vccd1 _06231_ sky130_fd_sc_hd__or4_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12006_ _04924_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17863_ _02122_ _02123_ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a21o_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19602_ rbzero.spi_registers.new_texadd\[1\]\[18\] rbzero.spi_registers.spi_buffer\[18\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
X_16814_ _09839_ _09840_ _09841_ vssd1 vssd1 vccd1 vccd1 _09842_ sky130_fd_sc_hd__a21oi_1
X_17794_ _01988_ _01989_ _02083_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19533_ _03394_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__clkbuf_1
X_16745_ _09782_ vssd1 vssd1 vccd1 vccd1 _09783_ sky130_fd_sc_hd__inv_2
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13957_ _07119_ _07126_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__or2_1
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19464_ rbzero.spi_registers.got_new_vshift _03118_ _03316_ _03351_ vssd1 vssd1 vccd1
+ vccd1 _00942_ sky130_fd_sc_hd__a31o_1
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12908_ rbzero.map_rom.a6 _06077_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__nand2_1
X_16676_ rbzero.row_render.size\[3\] _09746_ _09750_ _07954_ vssd1 vssd1 vccd1 vccd1
+ _00486_ sky130_fd_sc_hd__a22o_1
X_13888_ _06883_ _06882_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__or2b_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ _08718_ _08719_ _08720_ _08721_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__a2bb2o_1
X_18415_ _02569_ rbzero.debug_overlay.vplaneX\[-4\] _02642_ _02643_ vssd1 vssd1 vccd1
+ vccd1 _02645_ sky130_fd_sc_hd__nor4_1
X_12839_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and2_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ _02473_ rbzero.spi_registers.new_floor\[0\] _03319_ vssd1 vssd1 vccd1 vccd1
+ _03320_ sky130_fd_sc_hd__mux2_1
XFILLER_210_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ rbzero.wall_tracer.rayAddendX\[0\] _02580_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02581_ sky130_fd_sc_hd__mux2_1
X_15558_ _08632_ _08649_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__o21a_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20237__108 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__inv_2
X_14509_ _07306_ _07476_ _07444_ _06993_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__o22a_1
XFILLER_175_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18277_ _02514_ _02515_ _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__o21ba_1
X_15489_ _08575_ _08576_ _08583_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__a21o_1
X_17228_ _10246_ _10247_ vssd1 vssd1 vccd1 vccd1 _10248_ sky130_fd_sc_hd__and2_1
XFILLER_174_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput30 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_4
Xinput41 i_mode[1] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_16
Xinput52 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17159_ _10147_ _10178_ vssd1 vssd1 vccd1 vccd1 _10179_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03797_ clknet_0__03797_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03797_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20170_ _03751_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21624_ clknet_leaf_88_i_clk _01213_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21555_ clknet_leaf_13_i_clk _01144_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21486_ net204 _01075_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19658__39 clknet_1_0__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11170_ rbzero.tex_b0\[20\] rbzero.tex_b0\[19\] _04384_ vssd1 vssd1 vccd1 vccd1 _04387_
+ sky130_fd_sc_hd__mux2_1
X_20368_ clknet_1_0__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__buf_1
XFILLER_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22038_ clknet_leaf_35_i_clk _01627_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14860_ _06470_ _06575_ _07862_ _08014_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__a31o_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20342__203 clknet_1_0__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__inv_2
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13811_ _06658_ _06729_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__nand2_2
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14791_ _07955_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__clkbuf_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16530_ _09618_ _09619_ vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__xor2_1
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ _06765_ _06817_ _06818_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__or3b_1
XFILLER_1_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ rbzero.tex_b1\[58\] rbzero.tex_b1\[59\] _04270_ vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16461_ _09550_ _09551_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__and2_1
X_13673_ _06827_ _06829_ _06843_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__a21o_1
X_10885_ rbzero.tex_g0\[28\] rbzero.tex_g0\[27\] _04237_ vssd1 vssd1 vccd1 vccd1 _04238_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18200_ _02455_ _02465_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__and2_1
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15412_ _08195_ _08384_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__nor2_1
X_12624_ net19 net18 vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__or2_1
XFILLER_19_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19180_ rbzero.spi_registers.new_texadd\[1\]\[14\] _03188_ _03194_ _03184_ vssd1
+ vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__o211a_1
X_16392_ _09361_ _09382_ _09482_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__a21bo_1
XFILLER_200_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18131_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__or2_1
XFILLER_129_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15343_ _08437_ _08158_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__nor2_1
X_12555_ _04704_ _05732_ _05734_ _05703_ _05735_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__o2111a_1
X_20569__5 clknet_1_1__leaf__03457_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
XFILLER_200_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18062_ _09815_ _02346_ _02340_ rbzero.wall_tracer.trackDistY\[-10\] vssd1 vssd1
+ vccd1 vccd1 _00551_ sky130_fd_sc_hd__o2bb2a_1
X_11506_ _04653_ _04647_ _04695_ gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 _04696_
+ sky130_fd_sc_hd__o31a_1
X_15274_ _08246_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__buf_4
XFILLER_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ net51 _05637_ _05659_ net40 vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a22o_1
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17013_ _08952_ _09491_ vssd1 vssd1 vccd1 vccd1 _10034_ sky130_fd_sc_hd__nor2_1
XFILLER_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14225_ _07338_ _07337_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__and2_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ _04606_ _04613_ _04627_ _04628_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a211o_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14156_ _07211_ _07251_ _07326_ _07324_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__a31o_1
XFILLER_99_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11368_ rbzero.spi_registers.texadd2\[22\] rbzero.wall_hot\[0\] _04545_ rbzero.spi_registers.texadd1\[22\]
+ _04536_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a221o_1
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ rbzero.wall_tracer.mapY\[9\] _06078_ _06276_ vssd1 vssd1 vccd1 vccd1 _06279_
+ sky130_fd_sc_hd__o21a_1
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _03066_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__clkbuf_1
X_14087_ _07238_ _07240_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__and2b_1
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11299_ rbzero.spi_registers.texadd3\[7\] _04465_ _04455_ rbzero.spi_registers.texadd2\[7\]
+ _04469_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a221o_1
XFILLER_26_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17915_ _02201_ _02188_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__and2b_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13038_ _06166_ _06213_ _06163_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__or3b_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18895_ rbzero.pov.spi_buffer\[55\] rbzero.pov.ready_buffer\[55\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
XFILLER_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17846_ _08428_ _02012_ _02011_ _02008_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__o31ai_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17777_ _01955_ _01956_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nor2_1
X_14989_ _08104_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19516_ rbzero.spi_registers.new_texadd\[0\]\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__mux2_1
X_16728_ _06117_ _08218_ vssd1 vssd1 vccd1 vccd1 _09766_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19447_ _03348_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
X_16659_ _04415_ _04636_ _05283_ _03975_ vssd1 vssd1 vccd1 vccd1 _09740_ sky130_fd_sc_hd__a31o_1
XFILLER_23_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19378_ _02473_ rbzero.spi_registers.new_sky\[0\] _03309_ vssd1 vssd1 vccd1 vccd1
+ _03310_ sky130_fd_sc_hd__mux2_1
XFILLER_31_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18329_ _05120_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.debug_overlay.vplaneX\[-8\]
+ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__o31a_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21340_ clknet_leaf_22_i_clk _00929_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21271_ clknet_leaf_32_i_clk _00860_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20153_ _09734_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__buf_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20084_ rbzero.pov.ready_buffer\[16\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__and3_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20986_ clknet_leaf_26_i_clk _00575_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10670_ _04124_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21607_ clknet_leaf_15_i_clk _01196_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12340_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04907_ vssd1 vssd1 vccd1 vccd1 _05526_
+ sky130_fd_sc_hd__mux2_1
X_21538_ clknet_leaf_87_i_clk _01127_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ rbzero.row_render.side _05037_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand2_1
X_21469_ net187 _01058_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _07127_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__xor2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11222_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__buf_4
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ rbzero.tex_b0\[28\] rbzero.tex_b0\[27\] _04373_ vssd1 vssd1 vccd1 vccd1 _04378_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15961_ _09047_ _09055_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__xor2_2
X_11084_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _04340_ vssd1 vssd1 vccd1 vccd1 _04342_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17700_ _01917_ _01881_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__or2b_1
X_14912_ _08036_ _08053_ _08054_ _01633_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__o211a_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15892_ _08909_ _08938_ _08986_ _08901_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__a211oi_1
X_18680_ _02879_ _02880_ _02868_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__o21bai_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ rbzero.wall_tracer.visualWallDist\[3\] _08421_ vssd1 vssd1 vccd1 vccd1 _01922_
+ sky130_fd_sc_hd__nand2_2
X_14843_ rbzero.wall_tracer.stepDistY\[2\] _08000_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08001_ sky130_fd_sc_hd__mux2_1
XFILLER_36_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17562_ _01692_ _01741_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14774_ _07938_ _07939_ _07903_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11986_ _04645_ _05154_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a21o_1
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16513_ _09513_ _09484_ vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__or2b_1
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19301_ rbzero.spi_registers.texadd3\[18\] _03255_ vssd1 vssd1 vccd1 vccd1 _03264_
+ sky130_fd_sc_hd__or2_1
XFILLER_56_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13725_ _06810_ _06890_ _06894_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10937_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _04259_ vssd1 vssd1 vccd1 vccd1 _04265_
+ sky130_fd_sc_hd__mux2_1
X_17493_ _09647_ _09252_ _01679_ _01677_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__o31ai_2
XFILLER_32_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16444_ _08368_ _09397_ _09394_ _09534_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__o31a_1
X_19232_ rbzero.spi_registers.texadd2\[12\] _03222_ vssd1 vssd1 vccd1 vccd1 _03225_
+ sky130_fd_sc_hd__or2_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _06736_ _06740_ _06825_ _06826_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__a211o_1
X_10868_ rbzero.tex_g0\[36\] rbzero.tex_g0\[35\] _04226_ vssd1 vssd1 vccd1 vccd1 _04229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _05780_ _05781_ _05784_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
X_19163_ rbzero.spi_registers.texadd1\[7\] _03176_ vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__or2_1
X_16375_ _09355_ _09466_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__xor2_4
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13587_ _06725_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10799_ _04192_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__clkbuf_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18114_ _02390_ _02391_ _09869_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__o21ai_1
X_15326_ _08158_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19094_ rbzero.spi_registers.texadd0\[1\] _03143_ vssd1 vssd1 vccd1 vccd1 _03146_
+ sky130_fd_sc_hd__or2_1
X_12538_ net11 net10 vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nor2_2
XFILLER_173_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03803_ _03803_ vssd1 vssd1 vccd1 vccd1 clknet_0__03803_ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18045_ _02330_ _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__xnor2_1
X_15257_ _08350_ _08351_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__nor2_1
X_12469_ gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__buf_2
XFILLER_172_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _07365_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15188_ _08281_ _08282_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__and2_1
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20349__209 clknet_1_0__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__inv_2
XFILLER_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14139_ _07309_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__buf_2
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19996_ _03617_ _03637_ _06112_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a21o_1
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18947_ _03057_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18878_ rbzero.pov.spi_buffer\[47\] rbzero.pov.ready_buffer\[47\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
XFILLER_95_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17829_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__or2_1
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20840_ clknet_leaf_66_i_clk _00429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20771_ rbzero.wall_tracer.rayAddendY\[-7\] _02606_ _02557_ _03954_ vssd1 vssd1 vccd1
+ vccd1 _01653_ sky130_fd_sc_hd__a22o_1
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21323_ clknet_leaf_30_i_clk _00912_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21254_ clknet_leaf_0_i_clk _00843_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20205_ _03769_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21185_ clknet_leaf_18_i_clk _00774_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20289__156 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__inv_2
XFILLER_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20136_ _05650_ _03726_ _03727_ _03703_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__o211a_1
XFILLER_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ rbzero.pov.ready_buffer\[30\] _03684_ _03686_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01216_ sky130_fd_sc_hd__o211a_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ rbzero.row_render.wall\[1\] _05023_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_
+ sky130_fd_sc_hd__nand3_1
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _04959_ _04960_ _04944_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__mux2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ clknet_leaf_60_i_clk _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _06633_ _06675_ _06677_ _06678_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__a32o_4
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ rbzero.tex_g1\[40\] rbzero.tex_g1\[41\] _04144_ vssd1 vssd1 vccd1 vccd1 _04152_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14490_ _07651_ _07659_ _07660_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__a21boi_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20454__304 clknet_1_0__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__inv_2
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13441_ _06546_ _06579_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_1
X_10653_ _04115_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16160_ _08304_ _09252_ _09250_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ _06498_ _06501_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__nor2_1
X_10584_ _04079_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15111_ rbzero.wall_tracer.visualWallDist\[-7\] _08205_ _08168_ vssd1 vssd1 vccd1
+ vccd1 _08206_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12323_ _05507_ _05508_ _04934_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__mux2_1
XFILLER_10_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16091_ _08466_ _09184_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__and2_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15042_ _04464_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__buf_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ rbzero.tex_g1\[44\] _04905_ _05305_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1
+ _05441_ sky130_fd_sc_hd__a311o_1
XFILLER_170_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _04395_ vssd1 vssd1 vccd1 vccd1 _04405_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19850_ _03537_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
X_12185_ _05372_ _05036_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or2b_1
XFILLER_123_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18801_ rbzero.pov.spi_buffer\[10\] rbzero.pov.ready_buffer\[10\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02980_ sky130_fd_sc_hd__mux2_1
X_11136_ rbzero.tex_b0\[36\] rbzero.tex_b0\[35\] _04362_ vssd1 vssd1 vccd1 vccd1 _04369_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19781_ _03467_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__clkbuf_4
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16993_ _09882_ _09885_ _10012_ _10013_ vssd1 vssd1 vccd1 vccd1 _10015_ sky130_fd_sc_hd__o211a_1
XFILLER_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18732_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__and2b_1
X_15944_ _09036_ _09038_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__xnor2_2
X_11067_ rbzero.tex_b1\[4\] rbzero.tex_b1\[5\] _04325_ vssd1 vssd1 vccd1 vccd1 _04333_
+ sky130_fd_sc_hd__mux2_1
XFILLER_114_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15875_ _08943_ _08948_ _08968_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__nor3b_1
X_18663_ _02862_ _02863_ _02864_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__nand3_1
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _01895_ _01896_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a21oi_1
X_14826_ _07873_ _07985_ _06580_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__mux2_1
X_18594_ _05132_ rbzero.debug_overlay.vplaneY\[-8\] vssd1 vssd1 vccd1 vccd1 _02801_
+ sky130_fd_sc_hd__nand2_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _01831_ _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14757_ _07924_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__clkbuf_1
X_11969_ rbzero.debug_overlay.playerX\[-6\] _05121_ _05118_ rbzero.debug_overlay.playerX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a22o_1
X_13708_ _06770_ _06773_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__and3_1
X_17476_ _01670_ _01671_ _01668_ _01669_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__o2bb2a_1
X_14688_ _07837_ _07841_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__xnor2_1
X_19215_ rbzero.spi_registers.new_texadd\[2\]\[4\] _03206_ _03215_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00835_ sky130_fd_sc_hd__o211a_1
X_16427_ _09408_ _09516_ _09517_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__a21o_1
XFILLER_34_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ _06707_ _06807_ _06806_ _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__nand4_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ _09446_ _09448_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__nand2_1
X_19146_ rbzero.spi_registers.got_new_texadd\[1\] _03100_ vssd1 vssd1 vccd1 vccd1
+ _03175_ sky130_fd_sc_hd__and2_1
XFILLER_30_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ _08143_ _08401_ _08403_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__o21a_2
X_16289_ _09379_ _09380_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__xor2_1
XFILLER_195_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19077_ rbzero.map_overlay.i_mapdy\[5\] _03121_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or2_1
XFILLER_161_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18028_ _02007_ _09195_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__nor2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19979_ rbzero.pov.ready_buffer\[50\] _03438_ _03610_ _03626_ vssd1 vssd1 vccd1 vccd1
+ _03627_ sky130_fd_sc_hd__a211o_1
XFILLER_140_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21941_ net467 _01530_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21872_ net398 _01461_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20403__258 clknet_1_0__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__inv_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20823_ clknet_leaf_65_i_clk _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20754_ _02516_ _02515_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nor2_1
XFILLER_210_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20685_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _03903_
+ sky130_fd_sc_hd__nor2_1
XFILLER_195_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21306_ clknet_leaf_30_i_clk _00895_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21237_ clknet_leaf_4_i_clk _00826_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21168_ clknet_leaf_9_i_clk _00757_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20119_ _03440_ _03439_ _03445_ rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__a31o_1
X_13990_ _07154_ _07160_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__nand2_1
X_21099_ clknet_leaf_87_i_clk _00688_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__clkinv_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15660_ _08726_ _08753_ _08754_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__a21boi_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _06003_ _06046_ _06021_ _06006_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a311o_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _07773_ _07776_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__and2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _04909_ vssd1 vssd1 vccd1 vccd1 _05013_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _08671_ _08675_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__or2b_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _10220_ _10222_ vssd1 vssd1 vccd1 vccd1 _10349_ sky130_fd_sc_hd__nand2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _07674_ _07712_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__and2_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _04827_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__buf_6
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _10278_ _10279_ vssd1 vssd1 vccd1 vccd1 _10280_ sky130_fd_sc_hd__and2_1
X_10705_ _04142_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _07477_ _07641_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__and2b_1
XFILLER_201_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11685_ rbzero.row_render.size\[6\] _04418_ _04421_ rbzero.row_render.size\[5\] vssd1
+ vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__o2bb2a_1
X_16212_ _09302_ _09304_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__xor2_2
X_19000_ _03085_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__clkbuf_1
X_13424_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10636_ _04106_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__clkbuf_1
X_17192_ _10206_ _10211_ vssd1 vssd1 vccd1 vccd1 _10212_ sky130_fd_sc_hd__xnor2_1
X_16143_ _08148_ _09235_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__or3_2
X_13355_ _06517_ _06518_ _06520_ _06524_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__a41oi_2
X_10567_ _04070_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _05489_ _05490_ _05491_ _04946_ _04890_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__o221a_1
XFILLER_182_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ _09036_ _09038_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__nand2_1
XFILLER_143_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286_ _06449_ _06393_ _06406_ _06411_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__a31o_1
X_10498_ rbzero.tex_r1\[16\] rbzero.tex_r1\[17\] _04024_ vssd1 vssd1 vccd1 vccd1 _04032_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19902_ _03559_ _03567_ _03568_ _03302_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__o211a_1
X_15025_ _06106_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__buf_8
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ rbzero.tex_g1\[50\] _04829_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__or2_1
XFILLER_142_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19833_ _03528_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
X_12168_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04964_ vssd1 vssd1 vccd1 vccd1 _05356_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ rbzero.tex_b0\[44\] rbzero.tex_b0\[43\] _04351_ vssd1 vssd1 vccd1 vccd1 _04360_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19764_ _03492_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
X_16976_ _09896_ _09997_ vssd1 vssd1 vccd1 vccd1 _09998_ sky130_fd_sc_hd__nand2_1
X_12099_ _04655_ _05054_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__or2b_1
XFILLER_7_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18715_ rbzero.wall_tracer.rayAddendY\[8\] _02527_ _02906_ _02913_ vssd1 vssd1 vccd1
+ vccd1 _00637_ sky130_fd_sc_hd__o22a_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _08416_ _09002_ _09020_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__nand3_1
Xinput6 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18646_ _09753_ _02837_ _02838_ _02849_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__a31o_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _08471_ _08944_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__nand2_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ rbzero.wall_tracer.stepDistY\[-3\] _07971_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07972_ sky130_fd_sc_hd__mux2_1
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18577_ _02785_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__clkbuf_1
X_15789_ _08880_ _08883_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17528_ _01817_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__xor2_1
XFILLER_33_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17459_ _01750_ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__nand2_2
XFILLER_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19129_ rbzero.spi_registers.texadd0\[17\] _03156_ vssd1 vssd1 vccd1 vccd1 _03165_
+ sky130_fd_sc_hd__or2_1
XFILLER_145_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22071_ clknet_leaf_40_i_clk _01660_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21022_ clknet_leaf_74_i_clk _00611_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20483__330 clknet_1_0__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__inv_2
Xclkbuf_opt_2_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20327__189 clknet_1_1__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__inv_2
X_21924_ net450 _01513_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ net381 _01444_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20806_ clknet_leaf_50_i_clk _00395_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21786_ net312 _01375_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20737_ rbzero.traced_texVinit\[2\] _09759_ _03937_ _09101_ vssd1 vssd1 vccd1 vccd1
+ _01636_ sky130_fd_sc_hd__a22o_1
XFILLER_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _04645_ _04654_ _04655_ _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a41o_1
X_20668_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03889_
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ rbzero.tex_r1\[53\] rbzero.tex_r1\[54\] _03991_ vssd1 vssd1 vccd1 vccd1 _03992_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20599_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _03831_
+ sky130_fd_sc_hd__and2_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13140_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__and2_1
XFILLER_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20547__8 clknet_1_1__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _06239_ _06241_ _06243_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or4_1
XFILLER_133_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12022_ rbzero.tex_r1\[20\] _04906_ _05181_ _05209_ _05210_ vssd1 vssd1 vccd1 vccd1
+ _05211_ sky130_fd_sc_hd__a311o_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16830_ _09847_ _09850_ _09848_ vssd1 vssd1 vccd1 vccd1 _09856_ sky130_fd_sc_hd__o21ai_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13973_ _07112_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16761_ rbzero.wall_tracer.mapX\[9\] _09119_ vssd1 vssd1 vccd1 vccd1 _09796_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18500_ _02719_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__clkbuf_1
X_15712_ _08783_ _08805_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__nor2_1
X_12924_ rbzero.wall_tracer.mapY\[6\] _06077_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__xor2_1
X_19480_ rbzero.spi_registers.new_mapd\[4\] _02487_ _03362_ vssd1 vssd1 vccd1 vccd1
+ _03367_ sky130_fd_sc_hd__mux2_1
X_16692_ rbzero.row_render.texu\[4\] _09752_ _09754_ rbzero.texu_hot\[4\] vssd1 vssd1
+ vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18431_ _02651_ _02652_ _02659_ _08134_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15643_ _08668_ _08730_ _08737_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__nand3_1
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__nor2_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _04903_ _04987_ _04991_ _04995_ _04887_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o221a_1
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15574_ _08665_ _08668_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__nand2_1
X_18362_ _02557_ _02585_ _02586_ _02595_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a31o_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12786_ _04589_ _04704_ _04419_ _03973_ net34 net35 vssd1 vssd1 vccd1 vccd1 _05963_
+ sky130_fd_sc_hd__mux4_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17313_ _10330_ _10331_ _10218_ _10216_ vssd1 vssd1 vccd1 vccd1 _10332_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14525_ _07423_ _07204_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__nor2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__buf_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _02528_ _02529_ _02530_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17244_ _10261_ _10262_ _10135_ _10139_ vssd1 vssd1 vccd1 vccd1 _10263_ sky130_fd_sc_hd__o211a_1
X_14456_ _07625_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__and2_1
X_11668_ _04446_ _04837_ _04853_ _04854_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a311oi_1
XFILLER_186_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _06565_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__buf_4
X_10619_ _04097_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__clkbuf_1
X_17175_ _09397_ _09176_ _10066_ _10194_ vssd1 vssd1 vccd1 vccd1 _10195_ sky130_fd_sc_hd__o31a_1
XFILLER_174_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14387_ _07537_ _07557_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__and2_1
X_11599_ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__inv_2
X_16126_ _09217_ _09218_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__nand2_1
X_13338_ _06414_ _06386_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__nand2_1
XFILLER_182_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16057_ _08370_ _08325_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__or2_1
X_13269_ _06415_ _06438_ _06421_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ rbzero.wall_tracer.stepDistX\[9\] _08029_ _08091_ vssd1 vssd1 vccd1 vccd1
+ _08114_ sky130_fd_sc_hd__mux2_1
XFILLER_142_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19816_ _03519_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19747_ _03483_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
X_16959_ _09968_ _09980_ vssd1 vssd1 vccd1 vccd1 _09981_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18629_ _05127_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02833_
+ sky130_fd_sc_hd__and2_1
XFILLER_25_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21640_ clknet_leaf_85_i_clk _01229_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21571_ clknet_leaf_94_i_clk _01160_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 _08124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_22 rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20515__359 clknet_1_1__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__inv_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22054_ clknet_leaf_54_i_clk _01643_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21005_ clknet_leaf_25_i_clk _00594_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20409__264 clknet_1_1__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__inv_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _04282_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20260__129 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__inv_2
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21907_ net433 _01496_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _05771_ _05818_ _05819_ _05057_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__o22a_2
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21838_ net364 _01427_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _05744_ _05747_ _05748_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a22o_1
X_21769_ net295 _01358_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _07452_ _07480_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__nand2_1
XFILLER_106_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11522_ _04652_ rbzero.map_overlay.i_othery\[0\] vssd1 vssd1 vccd1 vccd1 _04712_
+ sky130_fd_sc_hd__xnor2_1
X_15290_ _08246_ _08384_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__nor2_1
XFILLER_183_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _07409_ _07411_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__nor2_1
X_11453_ net3 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__clkinv_4
XFILLER_183_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ rbzero.tex_r1\[61\] rbzero.tex_r1\[62\] _03980_ vssd1 vssd1 vccd1 vccd1 _03983_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14172_ _07342_ _07326_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11384_ _03971_ _04530_ _04533_ _04574_ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__o311a_1
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13123_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__nand2_1
XFILLER_139_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18980_ _03074_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17931_ _10315_ _09621_ _02218_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__or3_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13054_ _06120_ _06228_ _06129_ _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__or4_1
XFILLER_152_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12005_ rbzero.tex_r1\[8\] _04906_ _05181_ _05192_ _05193_ vssd1 vssd1 vccd1 vccd1
+ _05194_ sky130_fd_sc_hd__a311o_1
X_17862_ _02134_ _02150_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19601_ _03429_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16813_ _09832_ _09835_ _09833_ vssd1 vssd1 vccd1 vccd1 _09841_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17793_ _02081_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__or2_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19532_ rbzero.spi_registers.new_texadd\[0\]\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XFILLER_93_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16744_ _06264_ _09781_ vssd1 vssd1 vccd1 vccd1 _09782_ sky130_fd_sc_hd__and2_4
X_13956_ _07119_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nand2_1
XFILLER_59_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19463_ _03357_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ rbzero.map_rom.i_row\[4\] _06077_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__or2_1
X_13887_ _06930_ _07011_ _07055_ _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__a2bb2o_1
X_16675_ rbzero.row_render.size\[2\] _09746_ _09750_ _07944_ vssd1 vssd1 vccd1 vccd1
+ _00485_ sky130_fd_sc_hd__a22o_1
XFILLER_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18414_ _02569_ rbzero.debug_overlay.vplaneX\[-4\] _02642_ _02643_ vssd1 vssd1 vccd1
+ vccd1 _02644_ sky130_fd_sc_hd__o22a_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15626_ _08718_ _08719_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__xor2_1
X_12838_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__xor2_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__buf_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ _02573_ _02579_ _08134_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
X_15557_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__nand2_1
X_12769_ net35 vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__buf_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _07252_ _07444_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__or3_1
X_15488_ _08578_ _08579_ _08582_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__a21bo_1
X_18276_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__and2_1
XFILLER_175_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17227_ _10244_ _10245_ vssd1 vssd1 vccd1 vccd1 _10247_ sky130_fd_sc_hd__nand2_1
XFILLER_163_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput20 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_4
XFILLER_174_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
X_14439_ _06959_ _07366_ _07310_ _06808_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_175_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput42 i_mode[2] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_4
XFILLER_190_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 i_vec_csb vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_6
X_17158_ _10149_ _10177_ vssd1 vssd1 vccd1 vccd1 _10178_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03796_ clknet_0__03796_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03796_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16109_ _09183_ _09202_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__xnor2_2
XFILLER_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17089_ _10106_ _10108_ vssd1 vssd1 vccd1 vccd1 _10110_ sky130_fd_sc_hd__and2_1
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21623_ clknet_leaf_88_i_clk _01212_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21554_ clknet_leaf_13_i_clk _01143_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21485_ net203 _01074_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22037_ clknet_leaf_36_i_clk _01626_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _06757_ _06854_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__nand2_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14790_ rbzero.wall_tracer.stepDistY\[-5\] _07954_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07955_ sky130_fd_sc_hd__mux2_1
XFILLER_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13741_ _06765_ _06817_ _06818_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__o21bai_1
X_10953_ _04273_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16460_ _09406_ _09176_ _09549_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__o21ai_1
X_13672_ _06840_ _06842_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__xor2_1
X_10884_ _04214_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15411_ _08489_ _08498_ _08504_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__a21o_1
X_12623_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__nor2_1
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16391_ _09383_ _09359_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__or2b_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18130_ _09887_ _02405_ _02340_ rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1
+ vccd1 _00560_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15342_ rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__clkinv_2
XFILLER_169_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12554_ _04414_ _05719_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__nand2_1
XFILLER_200_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ _04642_ _04648_ _04645_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__or3_1
XFILLER_200_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15273_ _08178_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__buf_2
X_18061_ _02341_ _02344_ _02345_ _02337_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__o31a_1
XFILLER_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12485_ net49 _05664_ _05663_ net50 _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__a221o_1
X_17012_ _10030_ _10032_ vssd1 vssd1 vccd1 vccd1 _10033_ sky130_fd_sc_hd__and2b_1
X_14224_ _07357_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__nor2_1
XFILLER_184_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11436_ _04412_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__buf_4
XFILLER_125_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14155_ _07324_ _07325_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__nor2_1
XFILLER_99_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11367_ _04556_ _04558_ _03970_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a21o_1
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13106_ rbzero.wall_tracer.mapY\[9\] _06265_ _06266_ _06278_ vssd1 vssd1 vccd1 vccd1
+ _00389_ sky130_fd_sc_hd__a22o_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14086_ _07215_ _07244_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__nand2_1
XFILLER_4_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18963_ rbzero.spi_registers.spi_buffer\[12\] rbzero.spi_registers.spi_buffer\[11\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
X_11298_ rbzero.spi_registers.texadd1\[7\] _04460_ vssd1 vssd1 vccd1 vccd1 _04490_
+ sky130_fd_sc_hd__and2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _02188_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__and2b_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ rbzero.wall_tracer.trackDistY\[8\] _06165_ rbzero.wall_tracer.trackDistY\[7\]
+ _06167_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__o221a_1
XFILLER_191_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18894_ _03028_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17845_ _02132_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__xor2_1
XFILLER_67_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17776_ _02028_ _02065_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14988_ rbzero.wall_tracer.stepDistX\[-1\] _07982_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08104_ sky130_fd_sc_hd__mux2_1
XFILLER_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19515_ rbzero.spi_registers.got_new_texadd\[3\] _08117_ _03116_ _03385_ vssd1 vssd1
+ vccd1 vccd1 _00965_ sky130_fd_sc_hd__a31o_1
X_16727_ rbzero.map_rom.f1 _09118_ vssd1 vssd1 vccd1 vccd1 _09765_ sky130_fd_sc_hd__and2_1
X_13939_ _06879_ _07097_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__a21bo_1
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19446_ rbzero.spi_registers.spi_buffer\[10\] rbzero.spi_registers.new_other\[10\]
+ _03337_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__mux2_1
X_16658_ _03975_ _04415_ _04636_ _05283_ vssd1 vssd1 vccd1 vccd1 _09739_ sky130_fd_sc_hd__and4_1
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _08701_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xnor2_2
XFILLER_210_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19377_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__buf_2
X_16589_ _08950_ _09559_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__or2_1
XFILLER_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18328_ rbzero.debug_overlay.vplaneX\[-9\] vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__inv_2
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18259_ _02504_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_i_clk clknet_opt_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21270_ clknet_leaf_28_i_clk _00859_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03779_ clknet_0__03779_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03779_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20152_ _04657_ _05648_ _03099_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__and3_1
XFILLER_131_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _05111_ _03676_ _03694_ _03695_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a211o_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20985_ clknet_leaf_26_i_clk _00574_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21606_ clknet_leaf_15_i_clk _01195_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21537_ clknet_leaf_89_i_clk _01126_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12270_ _04810_ _05401_ _05419_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a31oi_4
XFILLER_107_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21468_ net186 _01057_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11221_ _04410_ _04416_ _04051_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o21ai_2
XFILLER_150_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21399_ clknet_leaf_6_i_clk _00988_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11152_ _04377_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15960_ _09048_ _09054_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__xor2_2
X_11083_ _04341_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20266__135 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__inv_2
X_14911_ rbzero.wall_tracer.visualWallDist\[-6\] _08047_ vssd1 vssd1 vccd1 vccd1 _08054_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15891_ _08916_ _08937_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__xnor2_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ _01837_ _01830_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__or2b_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14842_ _06655_ _07998_ _07999_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__a21o_4
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17561_ _01738_ _01740_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__nor2_1
XFILLER_90_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ _04659_ _05163_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or3b_1
X_14773_ _07806_ _07858_ _07876_ _06589_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__a211o_1
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19300_ rbzero.spi_registers.new_texadd\[3\]\[17\] _03254_ _03263_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__o211a_1
XFILLER_205_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ _09479_ _09592_ _09590_ vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f__03799_ clknet_0__03799_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03799_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10936_ _04264_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
X_13724_ _06810_ _06890_ _06894_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__and3_1
XFILLER_56_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17492_ _01782_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__xor2_1
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19231_ rbzero.spi_registers.new_texadd\[2\]\[11\] _03221_ _03224_ _03213_ vssd1
+ vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__o211a_1
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16443_ _09276_ _09393_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__nand2_1
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10867_ _04228_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
X_13655_ _06824_ _06822_ _06823_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__and3_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _05770_ _05785_ net17 vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__o21a_1
X_19162_ rbzero.spi_registers.new_texadd\[1\]\[6\] _03174_ _03183_ _03184_ vssd1 vssd1
+ vccd1 vccd1 _00813_ sky130_fd_sc_hd__o211a_1
X_16374_ _09340_ _09465_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__xor2_4
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _06658_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__buf_2
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10798_ rbzero.tex_g1\[4\] rbzero.tex_g1\[5\] _04188_ vssd1 vssd1 vccd1 vccd1 _04192_
+ sky130_fd_sc_hd__mux2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _02388_ _02389_ _09866_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a21o_1
X_15325_ rbzero.wall_tracer.stepDistX\[1\] vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__inv_2
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ _05714_ _05716_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__o21a_1
XFILLER_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19093_ rbzero.spi_registers.new_texadd\[0\]\[0\] _03141_ _03144_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00783_ sky130_fd_sc_hd__o211a_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03802_ _03802_ vssd1 vssd1 vccd1 vccd1 clknet_0__03802_ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__xnor2_1
X_15256_ _08342_ _08349_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__and2_1
X_12468_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14207_ _07318_ _07371_ _07372_ _07374_ _07377_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__a32o_1
X_11419_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__or2_1
X_15187_ rbzero.debug_overlay.playerY\[-3\] _08259_ vssd1 vssd1 vccd1 vccd1 _08282_
+ sky130_fd_sc_hd__nand2_1
X_12399_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _04893_ vssd1 vssd1 vccd1 vccd1 _05584_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14138_ _07254_ _07285_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__xor2_4
XFILLER_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19995_ rbzero.debug_overlay.playerY\[1\] _03611_ _03638_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01192_ sky130_fd_sc_hd__a211o_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14069_ _07182_ _07190_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__a21bo_1
X_18946_ _02487_ _02485_ _03052_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18877_ _03019_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17828_ _02095_ _02115_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__nor2_1
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17759_ _02047_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__and2_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20770_ _02750_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19429_ _03339_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21322_ clknet_leaf_30_i_clk _00911_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21253_ clknet_leaf_1_i_clk _00842_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20204_ rbzero.spi_registers.new_texadd\[3\]\[17\] rbzero.spi_registers.spi_buffer\[17\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__mux2_1
XFILLER_11_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21184_ clknet_leaf_18_i_clk _00773_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20135_ _05650_ _09729_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XFILLER_132_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ rbzero.debug_overlay.facingY\[-1\] _03685_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__or2_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _04914_ vssd1 vssd1 vccd1 vccd1 _04960_
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ clknet_leaf_59_i_clk _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10721_ _04151_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__clkbuf_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20899_ clknet_leaf_53_i_clk _00488_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _06606_ _06609_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__mux2_1
X_10652_ rbzero.tex_r0\[10\] rbzero.tex_r0\[9\] _04110_ vssd1 vssd1 vccd1 vccd1 _04115_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13371_ _06463_ _06507_ _06520_ _06541_ _06486_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__o32ai_4
X_10583_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _04077_ vssd1 vssd1 vccd1 vccd1 _04079_
+ sky130_fd_sc_hd__mux2_1
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _05009_ vssd1 vssd1 vccd1 vccd1 _05508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15110_ _08204_ rbzero.debug_overlay.playerY\[-7\] _06075_ vssd1 vssd1 vccd1 vccd1
+ _08205_ sky130_fd_sc_hd__mux2_1
XFILLER_139_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16090_ rbzero.wall_tracer.stepDistX\[4\] _08357_ vssd1 vssd1 vccd1 vccd1 _09184_
+ sky130_fd_sc_hd__nand2_4
X_15041_ _08125_ _08133_ _08137_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__o21a_1
XFILLER_181_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12253_ rbzero.tex_g1\[45\] _04904_ _04831_ _04939_ vssd1 vssd1 vccd1 vccd1 _05440_
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ _04404_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ _04890_ _04934_ _05002_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__or3_1
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18800_ _02979_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
X_11135_ _04368_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19780_ _03500_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
X_16992_ _10012_ _10013_ _09882_ _09885_ vssd1 vssd1 vccd1 vccd1 _10014_ sky130_fd_sc_hd__a211oi_1
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _02927_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
X_15943_ _08390_ _09037_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__nor2_1
X_11066_ _04332_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18662_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _02821_
+ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _08966_ _08967_ _08949_ _08968_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _01897_ _01903_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14825_ _07876_ _07877_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__or2_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _05132_ rbzero.debug_overlay.vplaneY\[-8\] vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__or2_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17544_ _01834_ _01835_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__xnor2_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ rbzero.wall_tracer.stepDistY\[-8\] _07923_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07924_ sky130_fd_sc_hd__mux2_1
XFILLER_205_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11968_ rbzero.debug_overlay.playerX\[4\] _05095_ _05108_ rbzero.debug_overlay.playerX\[-1\]
+ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a221o_1
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _06770_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__nand2_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10919_ _04255_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
X_17475_ _01691_ _10386_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__or2b_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14687_ _07847_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__xnor2_2
X_11899_ gpout0.hpos\[8\] _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__xor2_1
X_20320__184 clknet_1_1__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__inv_2
XFILLER_60_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19214_ rbzero.spi_registers.texadd2\[4\] _03208_ vssd1 vssd1 vccd1 vccd1 _03215_
+ sky130_fd_sc_hd__or2_1
X_16426_ _09409_ _09413_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__and2_1
XFILLER_60_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _06790_ _06617_ _06721_ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_201_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19145_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__clkbuf_4
X_16357_ _09446_ _09448_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__nor2_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ _06681_ _06725_ _06736_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__nand4_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _04463_ _06402_ _08147_ _08402_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__a211o_1
X_19076_ rbzero.spi_registers.new_mapd\[8\] _03119_ _03134_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00777_ sky130_fd_sc_hd__o211a_1
X_16288_ _09247_ _09259_ _09257_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__o21a_1
X_18027_ _02310_ _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__xnor2_1
X_15239_ _07907_ _08333_ _08143_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__mux2_1
XFILLER_172_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19978_ _08283_ _03570_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nor2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18929_ _03046_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21940_ net466 _01529_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21871_ net397 _01460_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20822_ clknet_leaf_65_i_clk _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20753_ rbzero.wall_tracer.rayAddendX\[-9\] _09746_ _03942_ vssd1 vssd1 vccd1 vccd1
+ _01647_ sky130_fd_sc_hd__a21o_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20684_ rbzero.texV\[6\] _03814_ _03819_ _03902_ vssd1 vssd1 vccd1 vccd1 _01617_
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20295__161 clknet_1_0__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__inv_2
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21305_ clknet_leaf_30_i_clk _00894_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21236_ clknet_leaf_5_i_clk _00825_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21167_ clknet_leaf_9_i_clk _00756_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20118_ rbzero.pov.ready_buffer\[10\] _03663_ _03713_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01240_ sky130_fd_sc_hd__o211a_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21098_ clknet_leaf_89_i_clk _00687_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20049_ rbzero.pov.ready_buffer\[23\] _03656_ _03675_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01209_ sky130_fd_sc_hd__o211a_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12940_ _06111_ rbzero.map_rom.c6 rbzero.map_rom.b6 _06112_ _06115_ vssd1 vssd1 vccd1
+ vccd1 _06116_ sky130_fd_sc_hd__a221o_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12871_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__or2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _07733_ _07735_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ rbzero.tex_r0\[63\] _04927_ _04929_ _04904_ vssd1 vssd1 vccd1 vccd1 _05012_
+ sky130_fd_sc_hd__a31o_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _08681_ _08682_ _08683_ _08684_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__a22o_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20378__236 clknet_1_1__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__inv_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _04909_ vssd1 vssd1 vccd1 vccd1 _04943_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14541_ _07709_ _07710_ _07711_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__nor3b_2
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ rbzero.tex_g1\[48\] rbzero.tex_g1\[49\] _04132_ vssd1 vssd1 vccd1 vccd1 _04142_
+ sky130_fd_sc_hd__mux2_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17260_ _09146_ _09490_ vssd1 vssd1 vccd1 vccd1 _10279_ sky130_fd_sc_hd__nor2_1
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14472_ _07601_ _07619_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__xnor2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ rbzero.row_render.size\[5\] _04421_ _04414_ rbzero.row_render.size\[4\] _04873_
+ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a221o_1
XFILLER_201_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16211_ _09290_ _09303_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__xor2_2
X_10635_ rbzero.tex_r0\[18\] rbzero.tex_r0\[17\] _04099_ vssd1 vssd1 vccd1 vccd1 _04106_
+ sky130_fd_sc_hd__mux2_1
X_13423_ _06566_ _06572_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nand2_2
X_17191_ _10209_ _10210_ vssd1 vssd1 vccd1 vccd1 _10211_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13354_ _06436_ _06445_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__nand2_4
X_16142_ _09121_ _09234_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__nor2_1
X_10566_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _04066_ vssd1 vssd1 vccd1 vccd1 _04070_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _04908_ vssd1 vssd1 vccd1 vccd1 _05491_
+ sky130_fd_sc_hd__mux2_1
X_16073_ _08434_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__clkbuf_4
X_13285_ _06336_ _06338_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__nand2_1
X_10497_ _04031_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12236_ rbzero.tex_g1\[52\] _04905_ _05305_ _05421_ _05422_ vssd1 vssd1 vccd1 vccd1
+ _05423_ sky130_fd_sc_hd__a311o_1
X_19901_ rbzero.debug_overlay.playerX\[-7\] _03565_ vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__or2_1
X_15024_ _08122_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19832_ rbzero.pov.spi_buffer\[53\] rbzero.pov.spi_buffer\[54\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
XFILLER_111_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12167_ _05353_ _05354_ _05191_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__mux2_1
XFILLER_2_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11118_ _04359_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19763_ rbzero.pov.spi_buffer\[20\] rbzero.pov.spi_buffer\[21\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
X_16975_ _09995_ _09996_ vssd1 vssd1 vccd1 vccd1 _09997_ sky130_fd_sc_hd__xor2_1
X_12098_ _04651_ _04578_ _05279_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a211o_1
XFILLER_7_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18714_ _08135_ _02911_ _02912_ _09745_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a31o_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15926_ _08416_ _09002_ _09020_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__a21o_1
X_11049_ _04323_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_6
XFILLER_7_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18645_ _08135_ _02847_ _02848_ _09751_ rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a32o_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08296_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__buf_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _07969_ _07970_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__or2_2
X_18576_ rbzero.wall_tracer.rayAddendY\[-2\] _02784_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15788_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__and2b_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17527_ _01818_ _09669_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__nor2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14739_ rbzero.wall_tracer.stepDistY\[-9\] _07907_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07908_ sky130_fd_sc_hd__mux2_1
XFILLER_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17458_ _10269_ _01749_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__or2_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16409_ _08847_ _08617_ _09076_ _08274_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__o22a_1
XFILLER_119_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _01675_ _01681_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19128_ rbzero.spi_registers.new_texadd\[0\]\[16\] _03155_ _03164_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__o211a_1
XFILLER_146_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19059_ rbzero.spi_registers.new_mapd\[12\] _03120_ _03125_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00769_ sky130_fd_sc_hd__o211a_1
XFILLER_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22070_ clknet_leaf_41_i_clk _01659_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21021_ clknet_leaf_74_i_clk _00610_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21923_ net449 _01512_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21854_ net380 _01443_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20805_ clknet_leaf_50_i_clk _00394_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21785_ net311 _01374_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20736_ rbzero.traced_texVinit\[1\] _09759_ _03937_ _09105_ vssd1 vssd1 vccd1 vccd1
+ _01635_ sky130_fd_sc_hd__a22o_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20667_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03888_
+ sky130_fd_sc_hd__or2_1
XFILLER_183_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _03979_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20598_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _03830_
+ sky130_fd_sc_hd__nor2_1
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ rbzero.map_overlay.i_otherx\[0\] _06108_ _06107_ rbzero.map_overlay.i_othery\[3\]
+ _06245_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a221o_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12021_ rbzero.tex_r1\[21\] _05185_ _05186_ _04937_ vssd1 vssd1 vccd1 vccd1 _05210_
+ sky130_fd_sc_hd__a31o_1
X_21219_ clknet_leaf_28_i_clk _00808_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16760_ rbzero.wall_tracer.mapX\[8\] _09119_ _09790_ _09793_ vssd1 vssd1 vccd1 vccd1
+ _09795_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13972_ _07130_ _07142_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__xor2_2
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15711_ _08783_ _08805_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__xor2_1
XFILLER_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _06081_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2_1
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16691_ rbzero.row_render.texu\[3\] _09752_ _09754_ rbzero.texu_hot\[3\] vssd1 vssd1
+ vccd1 vccd1 _00497_ sky130_fd_sc_hd__a22o_1
XFILLER_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18430_ _02657_ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15642_ _08732_ _08733_ _08735_ _08736_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__a31o_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nand2_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _04941_ _04994_ _04955_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a21o_1
X_18361_ _08135_ _02593_ _02594_ _09751_ rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a32o_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _08201_ _08439_ _08665_ _08667_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__or4bb_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _05650_ _05651_ _05958_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__mux2_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17312_ _09970_ _09972_ _08410_ _08390_ vssd1 vssd1 vccd1 vccd1 _10331_ sky130_fd_sc_hd__a211o_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__inv_2
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11736_ _04785_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18292_ _02528_ _02529_ _02530_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__or3_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17243_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _10262_ sky130_fd_sc_hd__nor2_1
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ _07531_ _07576_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__xor2_2
XFILLER_30_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ rbzero.row_render.size\[2\] gpout0.hpos\[2\] _04856_ vssd1 vssd1 vccd1 vccd1
+ _04857_ sky130_fd_sc_hd__a21oi_1
X_13406_ _06576_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__buf_4
X_10618_ rbzero.tex_r0\[26\] rbzero.tex_r0\[25\] _04088_ vssd1 vssd1 vccd1 vccd1 _04097_
+ sky130_fd_sc_hd__mux2_1
X_17174_ _09942_ _10065_ vssd1 vssd1 vccd1 vccd1 _10194_ sky130_fd_sc_hd__nand2_1
XFILLER_174_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11598_ _04772_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__or2_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14386_ _07533_ _07535_ _07536_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__a21o_1
XFILLER_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16125_ _09217_ _09218_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__nor2_1
X_10549_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _04055_ vssd1 vssd1 vccd1 vccd1 _04061_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__xor2_4
XFILLER_183_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20432__285 clknet_1_1__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__inv_2
X_16056_ _09148_ _09149_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13268_ _06415_ _06421_ _06438_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__and3_1
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15007_ _08113_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
X_12219_ rbzero.tex_g1\[18\] _05236_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__or2_1
X_13199_ rbzero.wall_tracer.rayAddendX\[-3\] _06369_ _06323_ vssd1 vssd1 vccd1 vccd1
+ _06370_ sky130_fd_sc_hd__mux2_2
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19815_ rbzero.pov.spi_buffer\[45\] rbzero.pov.spi_buffer\[46\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03519_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16958_ _09969_ _09979_ vssd1 vssd1 vccd1 vccd1 _09980_ sky130_fd_sc_hd__xor2_2
X_19746_ rbzero.pov.spi_buffer\[12\] rbzero.pov.spi_buffer\[13\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux2_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15909_ _08952_ _09003_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__or2_1
X_19677_ clknet_1_0__leaf__03457_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__buf_1
X_16889_ _09499_ _09630_ _09629_ vssd1 vssd1 vccd1 vccd1 _09911_ sky130_fd_sc_hd__a21bo_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18628_ rbzero.wall_tracer.rayAddendY\[2\] _02527_ _02825_ _02832_ vssd1 vssd1 vccd1
+ vccd1 _00631_ sky130_fd_sc_hd__o22a_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20221__94 clknet_1_1__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
X_18559_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__or2_1
XFILLER_75_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21570_ clknet_leaf_96_i_clk _01159_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _08136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_23 rbzero.wall_tracer.visualWallDist\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22053_ clknet_leaf_39_i_clk _01642_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21004_ clknet_leaf_3_i_clk _00593_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21906_ net432 _01495_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21837_ net363 _01426_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12570_ _04575_ _05732_ _05749_ _04628_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__o221a_1
X_21768_ net294 _01357_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ rbzero.map_overlay.i_otherx\[4\] _03972_ vssd1 vssd1 vccd1 vccd1 _04711_
+ sky130_fd_sc_hd__xnor2_1
X_20719_ _04429_ _04436_ rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a21boi_1
XFILLER_106_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21699_ net225 _01288_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ _07395_ _07410_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__nor2_1
X_11452_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__buf_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10403_ _03982_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14171_ _07211_ _07251_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__nand2_1
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11383_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__buf_4
XFILLER_165_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__and2_1
XFILLER_180_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19684__63 clknet_1_0__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XFILLER_140_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17930_ _02124_ _02216_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__o21ai_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _06144_ _06113_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__nand2_1
XFILLER_180_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ rbzero.tex_r1\[9\] _05185_ _05186_ _04953_ vssd1 vssd1 vccd1 vccd1 _05193_
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17861_ _02148_ _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__nor2_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19600_ rbzero.spi_registers.new_texadd\[1\]\[17\] rbzero.spi_registers.spi_buffer\[17\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
X_16812_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09840_ sky130_fd_sc_hd__nand2_1
XFILLER_4_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17792_ _01972_ _01980_ _02080_ _08123_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a31o_1
XFILLER_120_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19531_ _03393_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
X_16743_ _06217_ _06257_ _06161_ vssd1 vssd1 vccd1 vccd1 _09781_ sky130_fd_sc_hd__a21o_1
XFILLER_207_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _07122_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19462_ rbzero.spi_registers.new_vshift\[5\] _02489_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03357_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ rbzero.map_rom.i_row\[4\] _06077_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__nand2_1
XFILLER_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16674_ rbzero.row_render.size\[1\] _09746_ _09750_ _07935_ vssd1 vssd1 vccd1 vccd1
+ _00484_ sky130_fd_sc_hd__a22o_1
X_13886_ _06930_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18413_ _02596_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _02643_
+ sky130_fd_sc_hd__and2_1
XFILLER_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15625_ _08287_ _08343_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__nor2_1
XFILLER_50_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _06011_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nor2_1
X_19393_ _02474_ _04052_ _03307_ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1
+ vccd1 _03318_ sky130_fd_sc_hd__or4b_2
XFILLER_15_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18344_ _02576_ _02578_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15556_ _08364_ _08354_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__xnor2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12768_ net34 net35 vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__and2b_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ _07629_ _07675_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__a21o_1
X_11719_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__buf_6
X_18275_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nor2_1
X_15487_ _08580_ _08581_ _08502_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__or3_1
X_12699_ _05851_ _05854_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__nand2_1
X_17226_ _10244_ _10245_ vssd1 vssd1 vccd1 vccd1 _10246_ sky130_fd_sc_hd__or2_1
XFILLER_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput10 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_6
X_14438_ _07417_ _07248_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__nor2_1
Xinput21 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_4
XFILLER_200_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput32 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_4
XFILLER_122_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput43 i_reg_csb vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_8
Xinput54 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_4
X_17157_ _10159_ _10176_ vssd1 vssd1 vccd1 vccd1 _10177_ sky130_fd_sc_hd__xor2_1
XFILLER_190_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14369_ _07533_ _07537_ _07538_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_1__f__03795_ clknet_0__03795_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03795_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16108_ _09199_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__xnor2_2
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17088_ _10106_ _10108_ vssd1 vssd1 vccd1 vccd1 _10109_ sky130_fd_sc_hd__nor2_1
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16039_ _09130_ _09132_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19729_ rbzero.pov.spi_buffer\[4\] rbzero.pov.spi_buffer\[5\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03474_ sky130_fd_sc_hd__mux2_1
XFILLER_26_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21622_ clknet_leaf_87_i_clk _01211_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ clknet_leaf_94_i_clk _01142_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21484_ net202 _01073_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20435_ clknet_1_1__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__buf_1
XFILLER_180_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22036_ clknet_leaf_50_i_clk _01625_ vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13740_ _06907_ _06908_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__and3_1
X_10952_ rbzero.tex_b1\[59\] rbzero.tex_b1\[60\] _04270_ vssd1 vssd1 vccd1 vccd1 _04273_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _06797_ _06802_ _06841_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__o21a_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _04236_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
X_15410_ _08489_ _08498_ _08504_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__nand3_1
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ net17 _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__nor2_1
X_16390_ _09460_ _09357_ vssd1 vssd1 vccd1 vccd1 _09481_ sky130_fd_sc_hd__or2b_1
XFILLER_189_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15341_ _08433_ _08435_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12553_ _05702_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__or2_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18060_ _02342_ _02343_ _02334_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a21oi_1
X_11504_ _04691_ rbzero.debug_overlay.playerY\[-3\] _04692_ gpout0.hpos\[2\] _04693_
+ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o221a_1
X_15272_ _08172_ _08366_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__or2_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ net54 _05663_ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__and3_1
X_17011_ _09005_ _09242_ _10031_ vssd1 vssd1 vccd1 vccd1 _10032_ sky130_fd_sc_hd__or3_1
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14223_ _07358_ _07390_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__o21a_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ _04449_ _04616_ _04619_ _04626_ _04452_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__o311a_1
XFILLER_137_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11366_ rbzero.spi_registers.texadd1\[23\] _04545_ _04536_ _04557_ vssd1 vssd1 vccd1
+ vccd1 _04558_ sky130_fd_sc_hd__a211o_1
X_14154_ _07313_ _07320_ _07323_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__and3_1
XFILLER_4_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13105_ _06276_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14085_ _07213_ _07246_ _07255_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__a21oi_2
X_18962_ _03065_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__clkbuf_1
X_11297_ rbzero.texu_hot\[2\] _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17913_ _02193_ _02200_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__xnor2_1
X_13036_ rbzero.wall_tracer.trackDistY\[7\] _06167_ rbzero.wall_tracer.trackDistY\[6\]
+ _06168_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a221o_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18893_ rbzero.pov.spi_buffer\[54\] rbzero.pov.ready_buffer\[54\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17844_ _09647_ _09890_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__and2_1
XFILLER_26_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20544__386 clknet_1_0__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__inv_2
XFILLER_113_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17775_ _02063_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nor2_1
XFILLER_94_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14987_ _08091_ vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__buf_4
X_20243__114 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__inv_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19514_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__buf_4
X_16726_ _06126_ _09118_ vssd1 vssd1 vccd1 vccd1 _09764_ sky130_fd_sc_hd__xnor2_1
X_13938_ _07088_ _07096_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__or2b_1
XFILLER_170_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19445_ _03347_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ _09738_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__clkbuf_1
X_13869_ _07038_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__or2_1
XFILLER_179_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _08363_ _08702_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__nand2_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19376_ _04408_ _02930_ _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or3_2
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16588_ _08910_ _09677_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__nor2_1
XFILLER_194_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18327_ _02558_ _02559_ _02561_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a21o_1
XFILLER_37_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15539_ _08633_ _08589_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ rbzero.spi_registers.new_texadd\[2\]\[18\] rbzero.spi_registers.spi_buffer\[18\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17209_ _10101_ _10104_ vssd1 vssd1 vccd1 vccd1 _10229_ sky130_fd_sc_hd__and2b_1
XFILLER_175_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18189_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__nand2_1
X_19648__30 clknet_1_1__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03778_ clknet_0__03778_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03778_
+ sky130_fd_sc_hd__clkbuf_16
X_20151_ _05648_ _03099_ _03738_ _03703_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__o211a_1
X_19663__44 clknet_1_1__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_135_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20082_ _09734_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__buf_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ clknet_leaf_25_i_clk _00573_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21605_ clknet_leaf_13_i_clk _01194_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21536_ clknet_leaf_92_i_clk _01125_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21467_ net185 _01056_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11220_ _04411_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21398_ clknet_leaf_6_i_clk _00987_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _04373_ vssd1 vssd1 vccd1 vccd1 _04377_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11082_ rbzero.tex_b0\[62\] rbzero.tex_b0\[61\] _04340_ vssd1 vssd1 vccd1 vccd1 _04341_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22019_ clknet_leaf_50_i_clk _01608_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
X_14910_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.trackDistX\[-6\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__mux2_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _08984_ _08907_ _08938_ _08909_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__o22a_1
XFILLER_49_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14841_ _07826_ _07989_ _07887_ _06516_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__a31o_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _01804_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14772_ _07827_ _07872_ _07871_ _06577_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__a211o_1
X_11984_ rbzero.debug_overlay.playerY\[3\] _05098_ _05164_ _05172_ vssd1 vssd1 vccd1
+ vccd1 _05173_ sky130_fd_sc_hd__a211o_1
XFILLER_205_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03798_ clknet_0__03798_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03798_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16511_ _09477_ _09595_ _09596_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__o21ba_1
X_13723_ _06891_ _06892_ _06893_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__a21bo_1
X_17491_ _09525_ _09890_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__nand2_1
X_10935_ rbzero.tex_g0\[4\] rbzero.tex_g0\[3\] _04259_ vssd1 vssd1 vccd1 vccd1 _04264_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19230_ rbzero.spi_registers.texadd2\[11\] _03222_ vssd1 vssd1 vccd1 vccd1 _03224_
+ sky130_fd_sc_hd__or2_1
XFILLER_189_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _09531_ _09532_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ _06822_ _06823_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__a21oi_1
X_10866_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _04226_ vssd1 vssd1 vccd1 vccd1 _04228_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _05648_ _04657_ _05763_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__mux2_1
X_19161_ _03110_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__clkbuf_4
X_16373_ _09463_ _09464_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__or2_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _06754_ _06726_ _06727_ _06755_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__or4_1
X_10797_ _04191_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _02388_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__nor2_1
X_15324_ _08376_ _08418_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__xnor2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ _03110_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__clkbuf_4
X_12536_ net13 vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__inv_2
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03801_ _03801_ vssd1 vssd1 vccd1 vccd1 clknet_0__03801_ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18043_ _02177_ _02265_ _02266_ _02263_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a31o_1
X_15255_ _08342_ _08349_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__nor2_1
XFILLER_184_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _05648_ _04657_ _05646_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__mux2_1
X_14206_ _07375_ _07376_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11418_ rbzero.spi_registers.texadd3\[4\] _04457_ _04536_ rbzero.spi_registers.texadd0\[4\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a221o_1
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15186_ rbzero.debug_overlay.playerY\[-3\] _08259_ vssd1 vssd1 vccd1 vccd1 _08281_
+ sky130_fd_sc_hd__or2_1
X_12398_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _04931_ vssd1 vssd1 vccd1 vccd1 _05583_
+ sky130_fd_sc_hd__mux2_1
XFILLER_119_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14137_ _07305_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11349_ rbzero.spi_registers.texadd3\[19\] _04526_ _04537_ rbzero.spi_registers.texadd2\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a22o_1
X_19994_ rbzero.pov.ready_buffer\[54\] _03586_ _03636_ _03637_ _03617_ vssd1 vssd1
+ vccd1 vccd1 _03638_ sky130_fd_sc_hd__o221a_1
XFILLER_152_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14068_ _07184_ _07189_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__or2b_1
X_18945_ _03056_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ rbzero.wall_tracer.trackDistY\[-5\] _06183_ rbzero.wall_tracer.trackDistY\[-6\]
+ _06184_ _06194_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a221o_1
X_18876_ rbzero.pov.spi_buffer\[46\] rbzero.pov.ready_buffer\[46\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _02095_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__and2_1
XFILLER_67_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17758_ _09670_ _01922_ _02046_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__o21ai_1
XFILLER_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16709_ rbzero.traced_texa\[1\] _09757_ _09758_ rbzero.wall_tracer.visualWallDist\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
X_17689_ _01977_ _01978_ _01974_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a21o_1
XFILLER_74_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19428_ _02473_ rbzero.spi_registers.new_other\[0\] _03338_ vssd1 vssd1 vccd1 vccd1
+ _03339_ sky130_fd_sc_hd__mux2_1
XFILLER_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19359_ rbzero.spi_registers.got_new_vshift _03095_ vssd1 vssd1 vccd1 vccd1 _03298_
+ sky130_fd_sc_hd__and2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21321_ clknet_leaf_31_i_clk _00910_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_sky
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21252_ clknet_leaf_2_i_clk _00841_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20203_ _03768_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21183_ clknet_leaf_13_i_clk _00772_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20134_ _09729_ _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__and2_1
X_20065_ _03657_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__buf_2
XFILLER_58_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20527__370 clknet_1_1__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__inv_2
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ clknet_leaf_51_i_clk _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ rbzero.tex_g1\[41\] rbzero.tex_g1\[42\] _04144_ vssd1 vssd1 vccd1 vccd1 _04151_
+ sky130_fd_sc_hd__mux2_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ clknet_leaf_49_i_clk _00487_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_202_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ _04114_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ _04078_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__clkbuf_1
X_13370_ _06459_ _06507_ _06466_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__or3_2
XFILLER_16_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _05009_ vssd1 vssd1 vccd1 vccd1 _05507_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21519_ clknet_leaf_84_i_clk _01108_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20272__140 clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__inv_2
XFILLER_181_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15040_ _04526_ _08125_ _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12252_ rbzero.tex_g1\[47\] _04948_ _05438_ _04827_ vssd1 vssd1 vccd1 vccd1 _05439_
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ rbzero.tex_b0\[4\] rbzero.tex_b0\[3\] _04395_ vssd1 vssd1 vccd1 vccd1 _04404_
+ sky130_fd_sc_hd__mux2_1
X_12183_ _05027_ _05026_ rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1 vccd1 _05371_
+ sky130_fd_sc_hd__or3b_1
XFILLER_122_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _04362_ vssd1 vssd1 vccd1 vccd1 _04368_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16991_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _10013_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_82_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15942_ _08447_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__clkbuf_4
X_11065_ rbzero.tex_b1\[5\] rbzero.tex_b1\[6\] _04325_ vssd1 vssd1 vccd1 vccd1 _04332_
+ sky130_fd_sc_hd__mux2_1
X_18730_ rbzero.wall_tracer.rayAddendY\[10\] _02926_ _02524_ vssd1 vssd1 vccd1 vccd1
+ _02927_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18661_ _02838_ _02850_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__or2b_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _08956_ _08959_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__or2_1
XFILLER_37_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _01900_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__nand2_1
X_14824_ _07984_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _02797_ _02795_ _02796_ _04433_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_97_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ _09542_ _10215_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__nor2_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20555__16 clknet_1_0__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14755_ _07919_ _07922_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__nand2_2
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ rbzero.debug_overlay.playerX\[1\] _05096_ _05110_ rbzero.debug_overlay.playerX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a22o_1
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13706_ _06726_ _06719_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__nor2_1
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17474_ _01747_ _01748_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__or2_1
X_10918_ rbzero.tex_g0\[12\] rbzero.tex_g0\[11\] _04248_ vssd1 vssd1 vccd1 vccd1 _04255_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14686_ _07837_ _07841_ _07834_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_20_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _05066_ _05071_ _04640_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__o21bai_1
XFILLER_189_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16425_ _09409_ _09413_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__or2_1
X_19213_ rbzero.spi_registers.new_texadd\[2\]\[3\] _03206_ _03214_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00834_ sky130_fd_sc_hd__o211a_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13637_ _06771_ _06783_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__xnor2_4
X_10849_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _04215_ vssd1 vssd1 vccd1 vccd1 _04219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20355__215 clknet_1_1__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__inv_2
XFILLER_160_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19144_ rbzero.spi_registers.got_new_texadd\[1\] _03096_ vssd1 vssd1 vccd1 vccd1
+ _03173_ sky130_fd_sc_hd__nand2_2
X_16356_ _09301_ _09322_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13568_ _06737_ _06738_ _06735_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__a21o_1
XFILLER_34_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ rbzero.side_hot _06055_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__nor2_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12519_ reg_gpout\[0\] clknet_1_1__leaf__05700_ _05058_ vssd1 vssd1 vccd1 vccd1 _05701_
+ sky130_fd_sc_hd__mux2_2
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19075_ rbzero.map_overlay.i_mapdy\[4\] _03121_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__or2_1
X_16287_ _09368_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_35_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_121_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13499_ _06469_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nor2_2
XFILLER_201_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _02311_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__xor2_1
X_15238_ _06066_ _06375_ _04463_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ rbzero.wall_tracer.visualWallDist\[-4\] _08157_ _08263_ _08162_ vssd1 vssd1
+ vccd1 vccd1 _08264_ sky130_fd_sc_hd__a211o_1
XFILLER_5_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19977_ _03611_ _03624_ _03625_ _03579_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__o211a_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18928_ rbzero.pov.spi_buffer\[71\] rbzero.pov.ready_buffer\[71\] _02967_ vssd1 vssd1
+ vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18859_ rbzero.pov.spi_buffer\[38\] rbzero.pov.ready_buffer\[38\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
XFILLER_55_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21870_ net396 _01459_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20821_ clknet_leaf_65_i_clk _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20752_ _09749_ _02514_ _03941_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__and3_1
XFILLER_168_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20683_ _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21304_ clknet_leaf_30_i_clk _00893_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21235_ clknet_leaf_2_i_clk _00824_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21166_ clknet_leaf_95_i_clk _00755_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20117_ _02889_ _03655_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__nand2_1
X_21097_ clknet_leaf_89_i_clk _00686_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20048_ rbzero.debug_overlay.facingY\[-8\] _03658_ vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__or2_1
XFILLER_86_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _06010_ _06017_ _06005_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__nand3_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ rbzero.tex_r0\[62\] _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__and2_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ net145 _01588_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20304__169 clknet_1_0__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__inv_2
X_14540_ _07642_ _07668_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__xor2_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _04909_ vssd1 vssd1 vccd1 vccd1 _04942_
+ sky130_fd_sc_hd__mux2_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10703_ _04141_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__clkbuf_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _07641_ _07477_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__nor2b_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ rbzero.row_render.size\[3\] _04413_ _04414_ rbzero.row_render.size\[4\] _04872_
+ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__o221a_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _08466_ _09184_ _08390_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__a21oi_2
X_13422_ _06584_ _06586_ _06587_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__o31a_1
X_10634_ _04105_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__clkbuf_1
X_17190_ _09406_ _09669_ vssd1 vssd1 vccd1 vccd1 _10210_ sky130_fd_sc_hd__nor2_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16141_ _09121_ _09234_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__and2_1
X_13353_ _06502_ _06521_ _06522_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__or4_1
X_10565_ _04069_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ rbzero.tex_b0\[34\] _05314_ _04891_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a21o_1
XFILLER_143_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16072_ _08385_ _09027_ _09028_ _09030_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__a22o_1
X_13284_ _06452_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__xnor2_1
X_10496_ rbzero.tex_r1\[17\] rbzero.tex_r1\[18\] _04024_ vssd1 vssd1 vccd1 vccd1 _04031_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19900_ _08209_ rbzero.pov.ready_buffer\[61\] _03561_ vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__mux2_1
X_15023_ _08117_ _05632_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__and2_1
X_12235_ rbzero.tex_g1\[53\] _04904_ _05182_ _04939_ vssd1 vssd1 vccd1 vccd1 _05422_
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19831_ _03527_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12166_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _04964_ vssd1 vssd1 vccd1 vccd1 _05354_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _04351_ vssd1 vssd1 vccd1 vccd1 _04359_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19762_ _03491_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16974_ _09642_ _09710_ _09708_ vssd1 vssd1 vccd1 vccd1 _09996_ sky130_fd_sc_hd__a21oi_1
X_12097_ _04648_ _04418_ _05281_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or4_1
X_18713_ _02898_ _02900_ _02910_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__nand3_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15925_ _09010_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__xnor2_1
X_11048_ rbzero.tex_b1\[13\] rbzero.tex_b1\[14\] _04314_ vssd1 vssd1 vccd1 vccd1 _04323_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_6
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15856_ _08344_ _08950_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__nor2_1
X_18644_ _02839_ _02846_ _02840_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nand3_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14807_ _06581_ _07825_ _07866_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15787_ _08213_ _08195_ _08298_ _08337_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__or4_1
X_18575_ _02780_ _02781_ _02782_ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__inv_2
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17526_ _09397_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__buf_2
XFILLER_45_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _06525_ _07897_ _07906_ _06670_ _07891_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__a221o_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17457_ _10269_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__nand2_1
XFILLER_189_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__inv_2
XFILLER_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16408_ _08847_ _09076_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__nor2_1
X_17388_ _01679_ _01680_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__xor2_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16339_ _08441_ _09422_ _09427_ _09429_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__a2bb2o_1
X_19127_ rbzero.spi_registers.texadd0\[16\] _03156_ vssd1 vssd1 vccd1 vccd1 _03164_
+ sky130_fd_sc_hd__or2_1
XFILLER_158_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19058_ rbzero.map_overlay.i_mapdx\[2\] _03122_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or2_1
XFILLER_161_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18009_ _02277_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21020_ clknet_leaf_74_i_clk _00609_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21922_ net448 _01511_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21853_ net379 _01442_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20804_ clknet_leaf_51_i_clk _00393_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21784_ net310 _01373_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20735_ rbzero.traced_texVinit\[0\] _09759_ _03937_ _09111_ vssd1 vssd1 vccd1 vccd1
+ _01634_ sky130_fd_sc_hd__a22o_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20666_ _03734_ _03886_ _03887_ _03740_ rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1
+ _01614_ sky130_fd_sc_hd__a32o_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20597_ rbzero.texV\[-8\] _03695_ _03819_ _03829_ vssd1 vssd1 vccd1 vccd1 _01603_
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12020_ rbzero.tex_r1\[23\] _04933_ _05208_ _04923_ vssd1 vssd1 vccd1 vccd1 _05209_
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21218_ clknet_leaf_28_i_clk _00807_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21149_ clknet_leaf_100_i_clk _00738_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_20384__241 clknet_1_1__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__inv_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13971_ _07094_ _07141_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15710_ _08801_ _08803_ _08804_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__a21boi_1
XFILLER_4_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12922_ _06082_ _06083_ _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and3_1
XFILLER_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16690_ rbzero.row_render.texu\[2\] _09752_ _09754_ rbzero.texu_hot\[2\] vssd1 vssd1
+ vccd1 vccd1 _00496_ sky130_fd_sc_hd__a22o_1
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _08666_ _08734_ _08484_ _08471_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__and4bb_1
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12853_ _06018_ _06024_ _06025_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a211o_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _04992_ _04993_ _04912_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__mux2_1
X_18360_ _02577_ _02591_ _02587_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__or3_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15572_ _08382_ _08461_ _08457_ _08666_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__o22ai_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _05951_ _05957_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__a21o_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17311_ _09974_ _09975_ vssd1 vssd1 vccd1 vccd1 _10330_ sky130_fd_sc_hd__and2_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14523_ _07417_ _07209_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__nor2_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11735_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _04924_ vssd1 vssd1 vccd1 vccd1 _04925_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18291_ _02510_ _02521_ _02511_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__o21ai_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17242_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _10261_ sky130_fd_sc_hd__and2_1
X_14454_ _07580_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__nor2_1
XFILLER_175_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ gpout0.hpos\[1\] _03969_ _04836_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _06570_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__clkbuf_4
X_10617_ _04096_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__clkbuf_1
X_17173_ _10191_ _10192_ vssd1 vssd1 vccd1 vccd1 _10193_ sky130_fd_sc_hd__xnor2_1
X_14385_ _07541_ _07547_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__xor2_1
X_11597_ _04771_ _04768_ _04770_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and3_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _09072_ _09088_ _09071_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13336_ _06506_ _06413_ _06436_ _06445_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__or4bb_2
X_10548_ _04060_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16055_ _08952_ _08553_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__nor2_1
XFILLER_182_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _06416_ _06417_ _06418_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__or4_1
X_10479_ rbzero.tex_r1\[25\] rbzero.tex_r1\[26\] _04013_ vssd1 vssd1 vccd1 vccd1 _04022_
+ sky130_fd_sc_hd__mux2_1
X_20467__316 clknet_1_0__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__inv_2
XFILLER_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ rbzero.wall_tracer.stepDistX\[8\] _08027_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08113_ sky130_fd_sc_hd__mux2_1
X_12218_ rbzero.tex_g1\[20\] _05185_ _05181_ _05403_ _05404_ vssd1 vssd1 vccd1 vccd1
+ _05405_ sky130_fd_sc_hd__a311o_1
XFILLER_124_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13198_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__mux2_1
XFILLER_116_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19814_ _03518_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
X_12149_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _05010_ vssd1 vssd1 vccd1 vccd1 _05337_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19745_ _03482_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16957_ _09973_ _09976_ _09978_ vssd1 vssd1 vccd1 vccd1 _09979_ sky130_fd_sc_hd__mux2_1
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15908_ _08150_ _08165_ _08274_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__or3_1
X_16888_ _09908_ _09909_ vssd1 vssd1 vccd1 vccd1 _09910_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18627_ _02534_ _02831_ _09751_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__a21o_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15839_ _08916_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__nor2_1
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__and2_1
XFILLER_178_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ _01773_ _01774_ _01800_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a21o_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18489_ _06112_ _08124_ _02709_ _02710_ _02704_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__o221a_1
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _08136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_24 rbzero.wall_tracer.visualWallDist\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20333__195 clknet_1_0__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__inv_2
X_22052_ clknet_leaf_40_i_clk _01641_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21003_ clknet_leaf_3_i_clk _00592_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21905_ net431 _01494_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21836_ net362 _01425_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21767_ net293 _01356_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ _04670_ rbzero.map_overlay.i_othery\[4\] _04708_ _04578_ _04709_ vssd1 vssd1
+ vccd1 vccd1 _04710_ sky130_fd_sc_hd__o221a_1
XFILLER_141_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20718_ _04429_ _03928_ _03929_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__o21a_1
XFILLER_197_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21698_ net224 _01287_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ gpout0.hpos\[8\] _04640_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _04641_
+ sky130_fd_sc_hd__a21oi_2
X_20649_ _03870_ _03871_ _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a21o_1
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10402_ rbzero.tex_r1\[62\] rbzero.tex_r1\[63\] _03980_ vssd1 vssd1 vccd1 vccd1 _03982_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14170_ _07335_ _07340_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__xor2_1
X_11382_ _03971_ _04533_ _04573_ _04530_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__o22ai_1
XFILLER_180_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13121_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__or2_1
XFILLER_124_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__inv_2
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12003_ rbzero.tex_r1\[11\] _04933_ _05189_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17860_ _02146_ _02147_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__and2_1
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16811_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09839_ sky130_fd_sc_hd__or2_1
X_17791_ _01972_ _01980_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19530_ rbzero.spi_registers.new_texadd\[0\]\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _07123_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__nor2_1
X_16742_ _09778_ _09763_ _09777_ vssd1 vssd1 vccd1 vccd1 _09780_ sky130_fd_sc_hd__or3_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12905_ _06080_ _06077_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19461_ _03356_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16673_ rbzero.row_render.size\[0\] _09746_ _09750_ _07923_ vssd1 vssd1 vccd1 vccd1
+ _00483_ sky130_fd_sc_hd__a22o_1
X_13885_ _06971_ _07011_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nand2_1
XFILLER_59_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18412_ _02596_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _02642_
+ sky130_fd_sc_hd__nor2_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ _08265_ _08332_ _08335_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__or3_2
X_12836_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nor2_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ rbzero.spi_registers.got_new_sky _03118_ _03316_ _03317_ vssd1 vssd1 vccd1
+ vccd1 _00910_ sky130_fd_sc_hd__a31o_1
XFILLER_185_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15555_ _08632_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__xor2_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18343_ _05111_ rbzero.debug_overlay.vplaneX\[-9\] _02577_ vssd1 vssd1 vccd1 vccd1
+ _02578_ sky130_fd_sc_hd__a21oi_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ net35 net34 vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and2b_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ _07045_ _07209_ _07361_ _07253_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__o22a_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11718_ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__buf_6
X_18274_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__nand2_1
XFILLER_188_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15486_ rbzero.wall_tracer.visualWallDist\[-10\] _08156_ vssd1 vssd1 vccd1 vccd1
+ _08581_ sky130_fd_sc_hd__nand2_4
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ net27 _05860_ _05862_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a211o_2
X_17225_ _09894_ _10120_ _10118_ vssd1 vssd1 vccd1 vccd1 _10245_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14437_ _07561_ _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__nand2_1
Xinput11 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_6
X_11649_ rbzero.row_render.size\[5\] rbzero.row_render.size\[4\] _04838_ vssd1 vssd1
+ vccd1 vccd1 _04839_ sky130_fd_sc_hd__or3_1
Xinput22 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_168_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput33 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_4
X_17156_ _10174_ _10175_ vssd1 vssd1 vccd1 vccd1 _10176_ sky130_fd_sc_hd__nor2_1
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_8
XFILLER_196_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput55 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_6
X_14368_ _07533_ _07537_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03794_ clknet_0__03794_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03794_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16107_ _09047_ _09055_ _09200_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__a21bo_1
X_13319_ _06488_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nor2_1
X_17087_ _09954_ _09988_ _10107_ vssd1 vssd1 vccd1 vccd1 _10108_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14299_ _07467_ _07469_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__and2_1
XFILLER_171_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16038_ _08171_ _09131_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__nor2_1
XFILLER_157_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17989_ _02215_ _02240_ _02275_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19728_ _03473_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20521__365 clknet_1_0__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__inv_2
XFILLER_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21621_ clknet_leaf_87_i_clk _01210_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21552_ clknet_leaf_94_i_clk _01141_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21483_ net201 _01072_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20434_ clknet_1_1__leaf__04634_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__buf_1
XFILLER_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22035_ clknet_leaf_68_i_clk _01624_ vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _04272_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ _06788_ _06796_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__or2_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20496__342 clknet_1_1__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__inv_2
X_10882_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _04226_ vssd1 vssd1 vccd1 vccd1 _04236_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ net16 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__inv_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21819_ net345 _01408_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15340_ _08434_ _08409_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__nor2_1
XFILLER_12_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _04419_ _03973_ net10 vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__mux2_1
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11503_ rbzero.debug_overlay.playerX\[-2\] gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1
+ _04693_ sky130_fd_sc_hd__xnor2_1
X_15271_ _08303_ _08353_ _08365_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__a21boi_1
XFILLER_40_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12483_ net9 net8 vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__nor2_1
XFILLER_200_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17010_ _09146_ _09362_ vssd1 vssd1 vccd1 vccd1 _10031_ sky130_fd_sc_hd__or2_1
XFILLER_184_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14222_ _07391_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__or2b_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11434_ _04575_ _04622_ _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__or3_1
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14153_ _07313_ _07320_ _07323_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11365_ rbzero.spi_registers.texadd3\[23\] _04526_ _04537_ rbzero.spi_registers.texadd2\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a22o_1
XFILLER_4_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ rbzero.wall_tracer.mapY\[9\] _06078_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _07163_ _07198_ _07245_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__and3_1
X_18961_ rbzero.spi_registers.spi_buffer\[11\] rbzero.spi_registers.spi_buffer\[10\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11296_ rbzero.spi_registers.texadd0\[8\] _04466_ _04487_ vssd1 vssd1 vccd1 vccd1
+ _04488_ sky130_fd_sc_hd__o21a_1
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17912_ _02195_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__xor2_1
X_13035_ rbzero.wall_tracer.trackDistY\[6\] _06168_ _06169_ rbzero.wall_tracer.trackDistY\[5\]
+ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__o221a_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18892_ _03027_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17843_ _02129_ _02131_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__xor2_1
XFILLER_26_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17774_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__and2_1
X_14986_ _08102_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__clkbuf_1
X_19513_ _02477_ _03327_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__nor2_4
X_16725_ rbzero.map_rom.i_col\[4\] rbzero.wall_tracer.mapX\[5\] _09118_ vssd1 vssd1
+ vccd1 vccd1 _09763_ sky130_fd_sc_hd__o21a_1
X_13937_ _07058_ _07106_ _07107_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19444_ rbzero.spi_registers.spi_buffer\[9\] rbzero.spi_registers.new_other\[9\]
+ _03338_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__mux2_1
X_13868_ _07017_ _07037_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__xnor2_1
X_16656_ _05073_ _09732_ vssd1 vssd1 vccd1 vccd1 _09738_ sky130_fd_sc_hd__and2_1
XFILLER_62_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15607_ _08152_ _08616_ _08362_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__o21ai_2
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__and2_1
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19375_ _02475_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_done vssd1
+ vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or3b_1
X_16587_ _09422_ vssd1 vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__buf_2
X_13799_ _06924_ _06925_ _06919_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__o21ai_2
XFILLER_76_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18326_ _02558_ _02559_ _02561_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__nand3_1
XFILLER_187_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15538_ _08590_ _08584_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__and2b_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ _08561_ _08563_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__nor2_1
X_18257_ _02503_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ _10201_ _10227_ vssd1 vssd1 vccd1 vccd1 _10228_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__or2_1
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _10157_ _10158_ vssd1 vssd1 vccd1 vccd1 _10159_ sky130_fd_sc_hd__xor2_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03777_ clknet_0__03777_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03777_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20150_ _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__inv_2
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20081_ rbzero.pov.ready_buffer\[15\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03694_
+ sky130_fd_sc_hd__and3_1
XFILLER_83_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20445__296 clknet_1_1__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__inv_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20983_ clknet_leaf_25_i_clk _00572_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21604_ clknet_leaf_15_i_clk _01193_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_142_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21535_ clknet_leaf_93_i_clk _01124_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21466_ net184 _01055_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21397_ clknet_leaf_5_i_clk _00986_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11150_ _04376_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ _04214_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__clkbuf_4
X_20279_ clknet_1_1__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__buf_1
XFILLER_62_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22018_ clknet_leaf_48_i_clk _01607_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _07874_ _07881_ _06575_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__mux2_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14771_ _07914_ _07911_ _07894_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__mux2_1
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11983_ _05165_ _05166_ _05168_ _05171_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__or4_1
XFILLER_99_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03797_ clknet_0__03797_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03797_
+ sky130_fd_sc_hd__clkbuf_16
X_13722_ _06772_ _06790_ _06640_ _06733_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__or4_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16510_ _08148_ _09599_ _09600_ _08085_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__o211a_1
XFILLER_205_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10934_ _04263_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17490_ _01780_ _01781_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16441_ _09397_ _08384_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__nor2_1
X_13653_ _06799_ _06800_ _06801_ _06748_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__a22o_1
X_10865_ _04227_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _05782_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__or2_1
X_16372_ _09461_ _09462_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__and2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ rbzero.spi_registers.texadd1\[6\] _03176_ vssd1 vssd1 vccd1 vccd1 _03183_
+ sky130_fd_sc_hd__or2_1
X_13584_ _06708_ _06734_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nand2_2
X_10796_ rbzero.tex_g1\[5\] rbzero.tex_g1\[6\] _04188_ vssd1 vssd1 vccd1 vccd1 _04191_
+ sky130_fd_sc_hd__mux2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15323_ _08416_ _08417_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__nand2_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _02380_ _02382_ _02381_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a21boi_1
XFILLER_169_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12535_ net50 _05712_ _05715_ net49 vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a22o_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19091_ rbzero.spi_registers.texadd0\[0\] _03143_ vssd1 vssd1 vccd1 vccd1 _03144_
+ sky130_fd_sc_hd__or2_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03800_ _03800_ vssd1 vssd1 vccd1 vccd1 clknet_0__03800_ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ _08314_ _08327_ _08337_ _08348_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__o31a_1
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18042_ _08124_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__or3b_1
X_12466_ _04651_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__buf_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14205_ _06759_ _07310_ _07249_ _07306_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ rbzero.spi_registers.texadd2\[4\] _04537_ _04545_ rbzero.spi_registers.texadd1\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a22o_1
X_15185_ _08279_ rbzero.debug_overlay.playerX\[-3\] _08218_ vssd1 vssd1 vccd1 vccd1
+ _08280_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12397_ _04953_ _05577_ _05581_ _04967_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a211o_1
XFILLER_125_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14136_ _07306_ _07303_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11348_ rbzero.spi_registers.texadd0\[18\] _04535_ _04539_ vssd1 vssd1 vccd1 vccd1
+ _04540_ sky130_fd_sc_hd__o21a_1
X_19993_ rbzero.debug_overlay.playerY\[1\] _03632_ _03585_ vssd1 vssd1 vccd1 vccd1
+ _03637_ sky130_fd_sc_hd__o21ai_1
XFILLER_98_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _07236_ _07237_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__or2_1
X_18944_ _02485_ _02483_ _03052_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ rbzero.spi_registers.texadd3\[12\] _04465_ _04456_ rbzero.spi_registers.texadd2\[12\]
+ _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__a221o_1
XFILLER_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ rbzero.wall_tracer.trackDistY\[-6\] _06184_ _06185_ rbzero.wall_tracer.trackDistY\[-7\]
+ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__o221a_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18875_ _03018_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ _02097_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17757_ _09670_ _01922_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__or3_1
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14969_ rbzero.wall_tracer.stepDistX\[-10\] _07892_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08094_ sky130_fd_sc_hd__mux2_1
XFILLER_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16708_ _09749_ vssd1 vssd1 vccd1 vccd1 _09758_ sky130_fd_sc_hd__buf_2
XFILLER_39_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17688_ _01974_ _01977_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__and3_1
X_19427_ _03337_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__clkbuf_4
X_16639_ _04051_ _04637_ _05053_ _09727_ vssd1 vssd1 vccd1 vccd1 _09728_ sky130_fd_sc_hd__and4_1
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19358_ rbzero.spi_registers.got_new_vshift _03097_ vssd1 vssd1 vccd1 vccd1 _03297_
+ sky130_fd_sc_hd__nand2_2
XFILLER_188_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18309_ rbzero.wall_tracer.rayAddendX\[-3\] _02527_ _02543_ _02546_ vssd1 vssd1 vccd1
+ vccd1 _00598_ sky130_fd_sc_hd__o22a_1
XFILLER_176_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ rbzero.spi_registers.texadd3\[12\] _03255_ vssd1 vssd1 vccd1 vccd1 _03258_
+ sky130_fd_sc_hd__or2_1
XFILLER_198_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21320_ clknet_leaf_30_i_clk _00909_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21251_ clknet_leaf_24_i_clk _00840_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_20202_ rbzero.spi_registers.new_texadd\[3\]\[16\] rbzero.spi_registers.spi_buffer\[16\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21182_ clknet_leaf_13_i_clk _00771_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20133_ _05652_ _04695_ _03719_ _05653_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__or4b_1
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20064_ _03654_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ clknet_leaf_52_i_clk _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20897_ clknet_leaf_50_i_clk _00486_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _04110_ vssd1 vssd1 vccd1 vccd1 _04114_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ rbzero.tex_r0\[44\] rbzero.tex_r0\[43\] _04077_ vssd1 vssd1 vccd1 vccd1 _04078_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _04958_ _05480_ _05488_ _05505_ _04810_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a311o_1
XFILLER_16_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21518_ clknet_leaf_84_i_clk _01107_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12251_ rbzero.tex_g1\[46\] _04829_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or2_1
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21449_ net167 _01038_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11202_ _04403_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _05319_ _05336_ _05352_ _05369_ _05017_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__o221a_2
XFILLER_150_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ _04367_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16990_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _10012_ sky130_fd_sc_hd__or2_1
XFILLER_123_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15941_ _08910_ _08429_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__nor2_1
X_11064_ _04331_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18660_ _02860_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__nand2_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _08963_ _08965_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__or2_1
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _01787_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__or2_1
XFILLER_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ rbzero.wall_tracer.stepDistY\[-1\] _07982_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _07984_ sky130_fd_sc_hd__mux2_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _02795_ _02796_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__o21ai_1
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17542_ _01718_ _01832_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__o21ai_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11966_ rbzero.debug_overlay.playerX\[3\] _05098_ _05115_ rbzero.debug_overlay.playerX\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__a22o_1
X_14754_ _06655_ _07921_ _07891_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__a21oi_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10917_ _04254_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
X_13705_ _06851_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__xnor2_1
X_17473_ _01761_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__o21a_1
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14685_ _07827_ _07854_ _07855_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__o21a_1
X_11897_ gpout0.hpos\[4\] _05075_ _05083_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__or3_2
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19212_ rbzero.spi_registers.texadd2\[3\] _03208_ vssd1 vssd1 vccd1 vccd1 _03214_
+ sky130_fd_sc_hd__or2_1
X_16424_ _09392_ _09402_ _09400_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__a21o_1
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13636_ _06682_ _06784_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__and2_2
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10848_ _04218_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19143_ rbzero.spi_registers.new_texadd\[0\]\[23\] _03140_ _03172_ _03169_ vssd1
+ vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__o211a_1
X_16355_ _09319_ _09321_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__nor2_1
XFILLER_160_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13567_ _06721_ _06708_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__xnor2_4
X_10779_ rbzero.tex_g1\[13\] rbzero.tex_g1\[14\] _04177_ vssd1 vssd1 vccd1 vccd1 _04182_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19705__82 clknet_1_1__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
XFILLER_121_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ _07975_ _07982_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__xor2_1
X_12518_ net9 net8 _05382_ _05639_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o41a_2
X_16286_ _09376_ _09377_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__nand2_1
XFILLER_145_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19074_ rbzero.spi_registers.new_mapd\[7\] _03120_ _03133_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00776_ sky130_fd_sc_hd__o211a_1
XFILLER_160_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13498_ _06668_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18025_ _01697_ _09974_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__nor2_1
XFILLER_145_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ rbzero.wall_tracer.stepDistX\[-9\] _06262_ vssd1 vssd1 vccd1 vccd1 _08332_
+ sky130_fd_sc_hd__nor2_1
X_12449_ _05633_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15168_ _08258_ _06076_ _08262_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14119_ _06723_ _07268_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__and2_1
XFILLER_119_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19976_ _08258_ _03610_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__nand2_1
X_15099_ _08162_ _08187_ _08188_ _08193_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__a31o_1
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18927_ _03045_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _03009_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _01831_ _02032_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__nand2_1
X_18789_ _02973_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20820_ clknet_leaf_65_i_clk _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20751_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__or2_1
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20682_ _03893_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21303_ clknet_leaf_30_i_clk _00892_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21234_ clknet_leaf_2_i_clk _00823_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21165_ clknet_leaf_95_i_clk _00754_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ rbzero.pov.ready_buffer\[9\] _03663_ _03712_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01239_ sky130_fd_sc_hd__o211a_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21096_ clknet_leaf_89_i_clk _00685_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20047_ rbzero.debug_overlay.facingY\[-9\] _03663_ _03674_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01208_ sky130_fd_sc_hd__a211o_1
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _05009_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__buf_6
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ net144 _01587_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__buf_4
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20949_ clknet_leaf_59_i_clk _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ rbzero.tex_g1\[49\] rbzero.tex_g1\[50\] _04132_ vssd1 vssd1 vccd1 vccd1 _04141_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ _07592_ _07638_ _07640_ _07636_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__o31a_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ rbzero.row_render.size\[3\] _04413_ _04446_ rbzero.row_render.size\[2\] _04871_
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a221o_1
XFILLER_186_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20560__20 clknet_1_1__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
X_13421_ _06584_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__nand2_1
X_10633_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _04099_ vssd1 vssd1 vccd1 vccd1 _04105_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _09232_ _09233_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__nand2_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _06482_ _06513_ _06519_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__or3_1
X_10564_ rbzero.tex_r0\[52\] rbzero.tex_r0\[51\] _04066_ vssd1 vssd1 vccd1 vccd1 _04069_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ rbzero.tex_b0\[35\] _04926_ _04928_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__and3_1
X_16071_ _09144_ _09164_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ _06453_ _06393_ _06411_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21o_1
X_10495_ _04030_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ _08121_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
X_12234_ rbzero.tex_g1\[55\] _04948_ _05420_ _04827_ vssd1 vssd1 vccd1 vccd1 _05421_
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ rbzero.pov.spi_buffer\[52\] rbzero.pov.spi_buffer\[53\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12165_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _04932_ vssd1 vssd1 vccd1 vccd1 _05353_
+ sky130_fd_sc_hd__mux2_1
XFILLER_146_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ _04358_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19761_ rbzero.pov.spi_buffer\[19\] rbzero.pov.spi_buffer\[20\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16973_ _09929_ _09994_ vssd1 vssd1 vccd1 vccd1 _09995_ sky130_fd_sc_hd__xnor2_1
X_12096_ gpout0.vpos\[4\] _04578_ _04412_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1
+ _05285_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18712_ _02898_ _02900_ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a21o_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ _09017_ _09018_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__nor2_1
X_11047_ _04322_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_6
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20361__220 clknet_1_0__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__inv_2
X_18643_ _02839_ _02840_ _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a21o_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _08441_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__clkbuf_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14806_ _07903_ _07966_ _07968_ _07941_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__a211oi_2
XFILLER_18_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18574_ _05129_ _02773_ _04433_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__a21oi_1
X_15786_ _08195_ _08298_ _08337_ _08410_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__o22a_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _06173_ rbzero.wall_tracer.trackDistX\[-1\] vssd1 vssd1 vccd1 vccd1 _06174_
+ sky130_fd_sc_hd__nor2_1
XFILLER_206_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _01815_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__nand2_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737_ _06663_ _07898_ _07902_ _07903_ _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__o221a_1
X_11949_ rbzero.debug_overlay.facingY\[-6\] _05121_ _05118_ rbzero.debug_overlay.facingY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a22o_1
XFILLER_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17456_ _01747_ _01748_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__xor2_1
XFILLER_189_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ _07470_ _07527_ _07412_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__o21a_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _08952_ _09131_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__nor2_2
XFILLER_177_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13619_ _06783_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__clkbuf_4
X_17387_ _09647_ _09252_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__nor2_1
X_14599_ _07768_ _07769_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ rbzero.spi_registers.new_texadd\[0\]\[15\] _03155_ _03163_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__o211a_1
X_16338_ _08441_ _09422_ _09427_ _09429_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__or4bb_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19057_ rbzero.spi_registers.new_mapd\[11\] _03120_ _03124_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00768_ sky130_fd_sc_hd__o211a_1
X_16269_ _09270_ _09286_ _09360_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__a21bo_1
XFILLER_127_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _02278_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19959_ _08437_ _03611_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__nand2_1
XFILLER_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03459_ clknet_0__03459_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03459_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21921_ net447 _01510_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21852_ net378 _01441_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20803_ clknet_leaf_57_i_clk _00392_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21783_ net309 _01372_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20734_ _09749_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__buf_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_81_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20665_ _03882_ _03883_ _03884_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21o_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20596_ _03827_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21217_ clknet_leaf_6_i_clk _00806_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21148_ clknet_leaf_0_i_clk _00737_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21079_ clknet_leaf_85_i_clk _00668_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_13970_ _07139_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__nor2_1
XFILLER_86_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12921_ _06085_ _06095_ _06096_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__o21a_1
XFILLER_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_i_clk clknet_opt_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15640_ _08666_ _08472_ _08457_ _08734_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__o22ai_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _06026_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nand2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _04948_ vssd1 vssd1 vccd1 vccd1 _04993_
+ sky130_fd_sc_hd__mux2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _08177_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__clkbuf_4
X_12783_ net37 _05948_ _05959_ net38 vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a31o_1
XFILLER_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17310_ _10208_ _10210_ _10207_ vssd1 vssd1 vccd1 vccd1 _10329_ sky130_fd_sc_hd__a21bo_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11734_ _04914_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__buf_4
X_14522_ _07423_ _07248_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__nor3_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18290_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__and2_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17241_ _06172_ _09785_ _10260_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ _07598_ _07622_ _07623_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__a21oi_2
X_11665_ rbzero.row_render.size\[0\] gpout0.hpos\[1\] _04447_ rbzero.row_render.size\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__o211a_1
XFILLER_187_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10616_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _04088_ vssd1 vssd1 vccd1 vccd1 _04096_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13404_ _06574_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__buf_2
X_17172_ _08535_ _09037_ vssd1 vssd1 vccd1 vccd1 _10192_ sky130_fd_sc_hd__or2_1
XFILLER_174_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14384_ _07500_ _07512_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11596_ _04779_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nor2_2
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16123_ _09143_ _09216_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _06423_ _06446_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__xnor2_2
X_10547_ rbzero.tex_r0\[60\] rbzero.tex_r0\[59\] _04055_ vssd1 vssd1 vccd1 vccd1 _04060_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _09146_ _09003_ _09147_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13266_ _06329_ _06423_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__or2b_1
X_10478_ _04021_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12217_ rbzero.tex_g1\[21\] _04905_ _05186_ _04940_ vssd1 vssd1 vccd1 vccd1 _05404_
+ sky130_fd_sc_hd__a31o_1
X_15005_ _08112_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13197_ _06326_ _06065_ _06367_ _06323_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__o211a_1
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19813_ rbzero.pov.spi_buffer\[44\] rbzero.pov.spi_buffer\[45\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_1
X_12148_ _04958_ _05327_ _05335_ _04832_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__a31o_1
XFILLER_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19744_ rbzero.pov.spi_buffer\[11\] rbzero.pov.spi_buffer\[12\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16956_ _08637_ _09977_ _09691_ vssd1 vssd1 vccd1 vccd1 _09978_ sky130_fd_sc_hd__mux2_1
X_12079_ _04900_ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__and2b_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15907_ _08418_ _08376_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__or2b_1
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16887_ _08159_ _09608_ vssd1 vssd1 vccd1 vccd1 _09909_ sky130_fd_sc_hd__or2_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18626_ _02814_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__xnor2_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _08827_ _08915_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__and2_1
XFILLER_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18557_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__nor2_1
XFILLER_206_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15769_ _08812_ _08863_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__nor2_1
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _01784_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18488_ _08124_ _06094_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__nand2_1
XFILLER_75_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _01727_ _01730_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_14 _08136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_25 rbzero.wall_tracer.visualWallDist\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19109_ rbzero.spi_registers.new_texadd\[0\]\[8\] _03141_ _03153_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00791_ sky130_fd_sc_hd__o211a_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22051_ clknet_leaf_39_i_clk _01640_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21002_ clknet_leaf_3_i_clk _00591_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21904_ net430 _01493_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21835_ net361 _01424_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21766_ net292 _01355_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20717_ _04429_ _03928_ _08136_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21697_ net223 _01286_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11450_ gpout0.hpos\[7\] _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__and2_1
X_20648_ _03866_ _03868_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__nand2_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10401_ _03981_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__clkbuf_1
X_11381_ _03970_ _04525_ _04529_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__and3_1
X_20579_ _03734_ _03812_ _03813_ _03814_ rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1
+ _01600_ sky130_fd_sc_hd__a32o_1
XFILLER_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13120_ _06288_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nand3_1
XFILLER_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _06086_ _06107_ _06121_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__or3_1
XFILLER_180_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12002_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__buf_4
XFILLER_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16810_ _06185_ _09786_ _09838_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17790_ _02077_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__nand2_1
XFILLER_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16741_ _09763_ _09777_ _09778_ vssd1 vssd1 vccd1 vccd1 _09779_ sky130_fd_sc_hd__o21ai_1
X_13953_ _06748_ _06722_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__and2_1
XFILLER_115_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19460_ rbzero.spi_registers.new_vshift\[4\] _02487_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03356_ sky130_fd_sc_hd__mux2_1
X_12904_ rbzero.wall_tracer.mapY\[5\] vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__inv_2
X_16672_ rbzero.row_render.side _09746_ _09750_ _08138_ vssd1 vssd1 vccd1 vccd1 _00482_
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _07043_ _07053_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__a21o_1
X_18411_ _02638_ _02639_ _02637_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a21o_1
X_15623_ _08292_ _08357_ _08245_ _08296_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__a211o_1
XFILLER_59_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _03309_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__inv_2
XFILLER_188_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _05111_ _02555_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__nor2_1
XFILLER_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _08646_ _08647_ _08648_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__a21oi_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ _05941_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nand2_1
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20473__321 clknet_1_0__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__inv_2
X_14505_ _07629_ _07675_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nand2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _04892_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__buf_4
X_18273_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__nor2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15485_ _08161_ _08404_ _08406_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__o21a_2
X_12697_ _05864_ _05869_ _05875_ _05851_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a22o_2
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17224_ _10242_ _10243_ vssd1 vssd1 vccd1 vccd1 _10244_ sky130_fd_sc_hd__nand2_1
X_14436_ _06757_ _07303_ _07310_ _06807_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__a2bb2o_1
X_11648_ rbzero.row_render.size\[3\] _04837_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__or2_1
XFILLER_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_8
XFILLER_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_8
Xinput34 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_6
X_17155_ _10171_ _10173_ vssd1 vssd1 vccd1 vccd1 _10175_ sky130_fd_sc_hd__and2_1
Xinput45 i_reg_outs_enb vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_6
X_11579_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _04769_ sky130_fd_sc_hd__or2_1
XFILLER_122_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14367_ _07490_ _07493_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1__f__03793_ clknet_0__03793_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03793_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16106_ _09048_ _09054_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__nand2_1
X_13318_ _06459_ _06465_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__or2_1
X_17086_ _09985_ _09987_ vssd1 vssd1 vccd1 vccd1 _10107_ sky130_fd_sc_hd__and2b_1
X_14298_ _07395_ _07468_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__nor2_1
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ rbzero.wall_tracer.visualWallDist\[6\] _08475_ vssd1 vssd1 vccd1 vccd1 _09131_
+ sky130_fd_sc_hd__nand2_4
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ rbzero.wall_tracer.visualWallDist\[7\] _04428_ vssd1 vssd1 vccd1 vccd1 _06420_
+ sky130_fd_sc_hd__or2_1
XFILLER_111_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19690__68 clknet_1_1__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
XFILLER_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17988_ _02241_ _02213_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__and2b_1
XFILLER_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19727_ rbzero.pov.spi_buffer\[3\] rbzero.pov.spi_buffer\[4\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_78_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16939_ _09956_ _09960_ vssd1 vssd1 vccd1 vccd1 _09961_ sky130_fd_sc_hd__nand2_1
XFILLER_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__and2_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19589_ _03423_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21620_ clknet_leaf_87_i_clk _01209_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21551_ clknet_leaf_94_i_clk _01140_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21482_ net200 _01071_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22034_ clknet_leaf_67_i_clk _01623_ vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10950_ rbzero.tex_b1\[60\] rbzero.tex_b1\[61\] _04270_ vssd1 vssd1 vccd1 vccd1 _04272_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10881_ _04235_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _05711_ _05793_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a31o_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21818_ net344 _01407_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12551_ _05702_ net10 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__nand2_1
X_21749_ net275 _01338_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11502_ rbzero.debug_overlay.playerX\[-1\] vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__inv_2
X_15270_ _08354_ _08364_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__or2b_1
XFILLER_32_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ _05643_ _05646_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__nor2_1
XFILLER_138_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14221_ _07342_ _07364_ _07378_ _07379_ _07363_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__a32o_1
X_11433_ rbzero.spi_registers.texadd0\[3\] _04535_ _04623_ _04624_ _04454_ vssd1 vssd1
+ vccd1 vccd1 _04625_ sky130_fd_sc_hd__o221a_1
XFILLER_193_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14152_ _07321_ _07322_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__xnor2_1
X_11364_ rbzero.spi_registers.texadd0\[23\] _04535_ vssd1 vssd1 vccd1 vccd1 _04556_
+ sky130_fd_sc_hd__or2_1
XFILLER_164_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20316__180 clknet_1_0__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__inv_2
XFILLER_125_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13103_ _06272_ _06274_ _06270_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a21o_1
XFILLER_113_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14083_ _07212_ _07247_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__or2_2
XFILLER_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18960_ _03064_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11295_ rbzero.spi_registers.texadd1\[8\] _04460_ _04470_ _04486_ vssd1 vssd1 vccd1
+ vccd1 _04487_ sky130_fd_sc_hd__a211o_1
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17911_ _02197_ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__xnor2_1
X_13034_ _06169_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.trackDistY\[4\]
+ _06170_ _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a221o_1
XFILLER_65_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18891_ rbzero.pov.spi_buffer\[53\] rbzero.pov.ready_buffer\[53\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
XFILLER_117_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17842_ _09647_ _09621_ _01999_ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__o31a_1
XFILLER_154_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17773_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__nor2_1
X_14985_ rbzero.wall_tracer.stepDistX\[-2\] _07975_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08102_ sky130_fd_sc_hd__mux2_1
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19512_ rbzero.spi_registers.got_new_texadd\[2\] _08117_ _03316_ _02479_ vssd1 vssd1
+ vccd1 vccd1 _00964_ sky130_fd_sc_hd__a31o_1
X_16724_ _09762_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
X_13936_ _07104_ _06971_ _06930_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__or3_1
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19443_ _03346_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16655_ _09737_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__clkbuf_1
X_13867_ _06951_ _07033_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__nand2_1
XFILLER_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _08685_ _08690_ _08689_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__a21bo_1
X_12818_ _05994_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
X_19374_ _03306_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
X_16586_ _09664_ _09675_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__xor2_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13798_ _06967_ _06966_ _06968_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__nor3_2
XFILLER_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18325_ _02560_ _02550_ _02548_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a21o_1
XFILLER_76_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15537_ _08630_ _08631_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__or2_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ _05888_ _05881_ gpout4.clk_div\[1\] _05909_ _05926_ vssd1 vssd1 vccd1 vccd1
+ _05927_ sky130_fd_sc_hd__a41o_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18256_ rbzero.spi_registers.new_texadd\[2\]\[17\] rbzero.spi_registers.spi_buffer\[17\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15468_ _08298_ _08535_ _08531_ _08562_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__o31a_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17207_ _10224_ _10226_ vssd1 vssd1 vccd1 vccd1 _10227_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _07588_ _07589_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__nand2_1
X_18187_ _02454_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15399_ _08480_ _08493_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _08952_ _09890_ vssd1 vssd1 vccd1 vccd1 _10158_ sky130_fd_sc_hd__and2_1
XFILLER_183_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03776_ clknet_0__03776_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03776_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17069_ _10080_ _10089_ vssd1 vssd1 vccd1 vccd1 _10090_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20080_ rbzero.pov.ready_buffer\[14\] _03684_ _03693_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01222_ sky130_fd_sc_hd__o211a_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20982_ clknet_leaf_64_i_clk _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21603_ clknet_leaf_94_i_clk _01192_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21534_ clknet_leaf_93_i_clk _01123_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21465_ net183 _01054_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21396_ clknet_leaf_5_i_clk _00985_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ _04339_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22017_ clknet_leaf_48_i_clk _01606_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14770_ _07936_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__clkbuf_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ rbzero.debug_overlay.playerY\[-1\] _05108_ _05112_ rbzero.debug_overlay.playerY\[-5\]
+ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a221o_1
Xclkbuf_1_0__f__03796_ clknet_0__03796_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03796_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ _06707_ _06808_ _06805_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__a21o_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10933_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _04259_ vssd1 vssd1 vccd1 vccd1 _04263_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16440_ _09393_ _09529_ _09530_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__a21oi_1
X_10864_ rbzero.tex_g0\[38\] rbzero.tex_g0\[37\] _04226_ vssd1 vssd1 vccd1 vccd1 _04227_
+ sky130_fd_sc_hd__mux2_1
X_13652_ _06737_ _06725_ _06820_ _06821_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__a22o_1
XFILLER_72_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12603_ _05650_ _05651_ _05652_ _05653_ net16 net19 vssd1 vssd1 vccd1 vccd1 _05783_
+ sky130_fd_sc_hd__mux4_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _09461_ _09462_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__nor2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _04190_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__clkbuf_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13583_ _06633_ _06675_ _06677_ _06678_ _06680_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__a32oi_4
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _02386_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__or2b_1
X_15322_ _08415_ _08389_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__or2b_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _03142_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__buf_2
X_12534_ _05702_ _05704_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nor2_2
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _02169_ _02173_ _02255_ _02257_ _02326_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a311o_1
XFILLER_200_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15253_ _08345_ _08347_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nand2_1
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12465_ _04687_ _05644_ _05645_ _04642_ _05646_ _05640_ vssd1 vssd1 vccd1 vccd1 _05647_
+ sky130_fd_sc_hd__mux4_1
XFILLER_184_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_90 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_90/HI o_rgb[19] sky130_fd_sc_hd__conb_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ _07316_ _07204_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__or2_1
XFILLER_158_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11416_ rbzero.spi_registers.texadd3\[5\] _04457_ _04536_ rbzero.spi_registers.texadd0\[5\]
+ _03970_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a221o_1
X_12396_ _04922_ _05578_ _05579_ _05580_ _04940_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o221a_1
X_15184_ _08277_ _08278_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__and2_1
XFILLER_126_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14135_ _06727_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__buf_2
X_11347_ rbzero.spi_registers.texadd1\[18\] _04461_ _04536_ _04538_ vssd1 vssd1 vccd1
+ vccd1 _04539_ sky130_fd_sc_hd__a211o_1
XFILLER_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19992_ rbzero.debug_overlay.playerY\[1\] _03632_ vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__and2_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14066_ _07218_ _07192_ _07235_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__and3_1
X_11278_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__clkbuf_4
X_18943_ _03055_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13017_ _06185_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.trackDistY\[-8\]
+ _06186_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a221o_1
X_18874_ rbzero.pov.spi_buffer\[45\] rbzero.pov.ready_buffer\[45\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17825_ _02099_ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__xnor2_1
Xhold1 rbzero.tex_r1\[40\] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17756_ _01923_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a21o_1
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14968_ _08093_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16707_ rbzero.traced_texa\[0\] _09757_ _09756_ rbzero.wall_tracer.visualWallDist\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__a22o_1
XFILLER_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13919_ _06687_ _06719_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__nor2_1
X_17687_ _01865_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__o21ba_2
XFILLER_165_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14899_ _06103_ _08033_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__nor2_1
X_19426_ _04408_ _02932_ _03307_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__or3_1
X_16638_ _04414_ _04699_ vssd1 vssd1 vccd1 vccd1 _09727_ sky130_fd_sc_hd__nor2_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19357_ rbzero.color_floor\[5\] _03289_ _03296_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__a21o_1
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16569_ _09650_ _09658_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18308_ _02534_ _02544_ _02545_ _09745_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a31o_1
XFILLER_176_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19288_ rbzero.spi_registers.new_texadd\[3\]\[11\] _03254_ _03257_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__o211a_1
XFILLER_149_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18239_ _02478_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__buf_4
XFILLER_198_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21250_ clknet_leaf_24_i_clk _00839_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20201_ _03767_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21181_ clknet_leaf_13_i_clk _00770_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20132_ _03724_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20063_ rbzero.debug_overlay.facingY\[-2\] _03676_ _03683_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01215_ sky130_fd_sc_hd__a211o_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ clknet_leaf_52_i_clk _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ clknet_leaf_49_i_clk _00485_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10580_ _04054_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21517_ clknet_leaf_84_i_clk _01106_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _04967_ _05423_ _05427_ _04887_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a311o_1
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21448_ net166 _01037_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04395_ vssd1 vssd1 vccd1 vccd1 _04403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12181_ _04958_ _05360_ _05368_ _04810_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a31o_1
X_21379_ clknet_leaf_29_i_clk _00968_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11132_ rbzero.tex_b0\[38\] rbzero.tex_b0\[37\] _04362_ vssd1 vssd1 vccd1 vccd1 _04367_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15940_ _09033_ _09034_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__and2_1
X_11063_ rbzero.tex_b1\[6\] rbzero.tex_b1\[7\] _04325_ vssd1 vssd1 vccd1 vccd1 _04331_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _08963_ _08965_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20428__281 clknet_1_0__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__inv_2
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ rbzero.wall_tracer.visualWallDist\[5\] _01699_ vssd1 vssd1 vccd1 vccd1 _01901_
+ sky130_fd_sc_hd__nand2_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14822_ _07868_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__buf_4
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _02786_ _02788_ _02787_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__a21bo_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _08889_ _10093_ _10330_ _08816_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__o22ai_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _06574_ _07920_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__nor2_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11965_ _05064_ _05145_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o21ai_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03779_ clknet_0__03779_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03779_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13704_ _06865_ _06874_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__xnor2_2
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10916_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _04248_ vssd1 vssd1 vccd1 vccd1 _04254_
+ sky130_fd_sc_hd__mux2_1
X_17472_ _01761_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nor3_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14684_ _06613_ _07850_ _07853_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__nand3_2
X_11896_ _04578_ _05075_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nand3_2
XFILLER_189_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19211_ rbzero.spi_registers.new_texadd\[2\]\[2\] _03206_ _03211_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00833_ sky130_fd_sc_hd__o211a_1
X_16423_ _09484_ _09513_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__xnor2_1
X_13635_ _06617_ _06792_ _06805_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__or3b_1
X_10847_ rbzero.tex_g0\[46\] rbzero.tex_g0\[45\] _04215_ vssd1 vssd1 vccd1 vccd1 _04218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19142_ rbzero.spi_registers.texadd0\[23\] _03142_ vssd1 vssd1 vccd1 vccd1 _03172_
+ sky130_fd_sc_hd__or2_1
XFILLER_73_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16354_ _09444_ _09445_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__or2_1
XFILLER_201_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _06692_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__clkinv_2
X_10778_ _04181_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15305_ _08391_ _08399_ _06263_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__mux2_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19073_ rbzero.map_overlay.i_mapdy\[3\] _03122_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__or2_1
X_12517_ net9 _05677_ _05692_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__a211o_2
X_16285_ _09271_ _09369_ _09375_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__nand3_1
XFILLER_185_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13497_ _06537_ _06539_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__and2_1
X_18024_ _10288_ _10214_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__nor2_1
X_15236_ _08326_ _08330_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__nand2_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ reg_rgb\[23\] _05632_ _05058_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__mux2_4
XFILLER_201_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15167_ _06034_ _06074_ _08261_ _08156_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__a31o_1
X_12379_ _04922_ _05561_ _05563_ _04919_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o211a_1
XFILLER_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _06540_ _07078_ _07219_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__or3_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19975_ _08261_ rbzero.pov.ready_buffer\[49\] _03561_ vssd1 vssd1 vccd1 vccd1 _03624_
+ sky130_fd_sc_hd__mux2_1
X_15098_ _08191_ _08192_ _08156_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__mux2_1
XFILLER_87_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18926_ rbzero.pov.spi_buffer\[70\] rbzero.pov.ready_buffer\[70\] _02967_ vssd1 vssd1
+ vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
X_14049_ _06759_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__nand2_1
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18857_ rbzero.pov.spi_buffer\[37\] rbzero.pov.ready_buffer\[37\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03009_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17808_ _02054_ _02056_ _02096_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18788_ rbzero.pov.spi_buffer\[4\] rbzero.pov.ready_buffer\[4\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _09542_ _01943_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__or2_1
X_20750_ _03940_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ rbzero.spi_registers.spi_cmd\[0\] _02474_ vssd1 vssd1 vccd1 vccd1 _03327_
+ sky130_fd_sc_hd__or2b_1
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20681_ _03898_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nand2_1
XFILLER_51_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20256__126 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__inv_2
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21302_ clknet_leaf_36_i_clk _00891_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21233_ clknet_leaf_1_i_clk _00822_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21164_ clknet_leaf_95_i_clk _00753_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20115_ _02907_ _03655_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XFILLER_172_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21095_ clknet_leaf_92_i_clk _00684_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20046_ rbzero.pov.ready_buffer\[22\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__and3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ net143 _01586_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11750_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__buf_6
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20948_ clknet_leaf_59_i_clk _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ _04140_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11681_ rbzero.row_render.size\[0\] _04453_ _04869_ _04870_ vssd1 vssd1 vccd1 vccd1
+ _04871_ sky130_fd_sc_hd__o31a_1
XFILLER_144_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20879_ clknet_leaf_41_i_clk _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_13420_ _06588_ _06589_ _06590_ _06477_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__o22a_1
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ _04104_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10563_ _04068_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__clkbuf_1
X_13351_ _06488_ _06489_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__or2_1
XFILLER_195_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _04937_ _05483_ _05487_ _04902_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a211o_1
X_16070_ _09162_ _09163_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__nand2_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10494_ rbzero.tex_r1\[18\] rbzero.tex_r1\[19\] _04024_ vssd1 vssd1 vccd1 vccd1 _04030_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _04444_ _06402_ _06404_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a21o_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _08117_ _05551_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__and2_1
XFILLER_154_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ rbzero.tex_g1\[54\] _04830_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__or2_1
XFILLER_155_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ _04903_ _05343_ _05347_ _05351_ _04887_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__o221a_1
XFILLER_155_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11115_ rbzero.tex_b0\[46\] rbzero.tex_b0\[45\] _04351_ vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16972_ _09992_ _09993_ vssd1 vssd1 vccd1 vccd1 _09994_ sky130_fd_sc_hd__and2_1
XFILLER_190_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19760_ _03467_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__clkbuf_4
X_12095_ _04415_ _05283_ _04700_ _03972_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15923_ _09014_ _09016_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__and2_1
X_11046_ rbzero.tex_b1\[14\] rbzero.tex_b1\[15\] _04314_ vssd1 vssd1 vccd1 vccd1 _04322_
+ sky130_fd_sc_hd__mux2_1
X_18711_ _02907_ _02895_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a21oi_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20218__91 clknet_1_1__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18642_ _02844_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nand2_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _08943_ _08948_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__nand2_1
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _07903_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__nor2_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _05129_ _02773_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or2_1
X_15785_ _08228_ _08344_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__or2_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12997_ rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__inv_2
XFILLER_91_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _09528_ _09677_ _09560_ _08814_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__o22ai_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _06665_ _07904_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__or2_1
XFILLER_206_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11948_ rbzero.debug_overlay.facingY\[-3\] _05110_ _05108_ rbzero.debug_overlay.facingY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a22o_1
XFILLER_206_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _10358_ _10359_ _10361_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__o21a_1
XFILLER_162_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14667_ _07471_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__inv_2
X_11879_ _04638_ _04699_ _04639_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__o21ba_1
X_16406_ _09370_ _09371_ _09373_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ _06640_ _06785_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__nor2_1
X_17386_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nand2_1
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _07253_ _07476_ _07444_ _07045_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__o22a_1
XFILLER_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19125_ rbzero.spi_registers.texadd0\[15\] _03156_ vssd1 vssd1 vccd1 vccd1 _03163_
+ sky130_fd_sc_hd__or2_1
X_16337_ _08484_ _09426_ _09428_ vssd1 vssd1 vccd1 vccd1 _09429_ sky130_fd_sc_hd__a21o_1
XFILLER_185_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _06719_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__buf_2
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19056_ rbzero.map_overlay.i_mapdx\[1\] _03122_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__or2_1
X_16268_ _09287_ _09268_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__or2b_1
XFILLER_173_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18007_ _02279_ _02293_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__xnor2_1
X_15219_ _08298_ _08313_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__or2_1
XFILLER_160_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16199_ _09291_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__inv_2
XFILLER_142_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19958_ _08437_ rbzero.pov.ready_buffer\[44\] _03561_ vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18909_ _03036_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03458_ clknet_0__03458_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03458_
+ sky130_fd_sc_hd__clkbuf_16
X_19889_ net40 _03557_ _03095_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__o21ai_4
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21920_ net446 _01509_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21851_ net377 _01440_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20802_ clknet_leaf_58_i_clk _00391_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21782_ net308 _01371_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20733_ rbzero.hsync net63 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__nor2_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20664_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__inv_2
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20595_ _03820_ _03821_ _03822_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o21ai_1
XFILLER_167_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19696__74 clknet_1_1__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21216_ clknet_leaf_6_i_clk _00805_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21147_ clknet_leaf_99_i_clk _00736_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20310__175 clknet_1_1__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__inv_2
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21078_ clknet_leaf_83_i_clk _00667_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20029_ _03557_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__buf_2
X_12920_ rbzero.map_rom.a6 _06077_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__or2_1
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12851_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__or2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _04948_ vssd1 vssd1 vccd1 vccd1 _04992_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15570_ _08177_ _08382_ _08461_ _08457_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__or4_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _03969_ _04575_ _04452_ _04628_ _05958_ _05946_ vssd1 vssd1 vccd1 vccd1 _05959_
+ sky130_fd_sc_hd__mux4_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ _06959_ _07204_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__or2_1
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__buf_4
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _06105_ _10140_ _10259_ _09812_ vssd1 vssd1 vccd1 vccd1 _10260_ sky130_fd_sc_hd__o211a_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _07599_ _07621_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__nor2_1
X_20239__110 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__inv_2
X_11664_ _04412_ _04852_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__nor2_1
XFILLER_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13403_ _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__buf_2
X_10615_ _04095_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__clkbuf_1
X_17171_ _10189_ _10190_ vssd1 vssd1 vccd1 vccd1 _10191_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20391__247 clknet_1_1__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__inv_2
XFILLER_31_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14383_ _07551_ _07553_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__nor2_1
X_11595_ _04781_ _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__or2_4
XFILLER_128_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16122_ _09214_ _09215_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__nor2_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ _06495_ _06502_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__or3_2
X_10546_ _04059_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16053_ _08152_ _08847_ _09005_ _08166_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__o22ai_1
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265_ _06430_ _06432_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__a21oi_4
X_10477_ rbzero.tex_r1\[26\] rbzero.tex_r1\[27\] _04013_ vssd1 vssd1 vccd1 vccd1 _04021_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15004_ rbzero.wall_tracer.stepDistX\[7\] _08023_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08112_ sky130_fd_sc_hd__mux2_1
XFILLER_170_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12216_ rbzero.tex_g1\[23\] _04910_ _05402_ _04912_ vssd1 vssd1 vccd1 vccd1 _05403_
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13196_ rbzero.wall_tracer.visualWallDist\[-8\] rbzero.wall_tracer.rcp_sel\[2\] vssd1
+ vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__or2_1
XFILLER_155_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19812_ _03517_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
X_12147_ _04941_ _05330_ _05334_ _04902_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a211o_1
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19743_ _03481_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
X_16955_ _08042_ _08338_ _09689_ vssd1 vssd1 vccd1 vccd1 _09977_ sky130_fd_sc_hd__or3_1
X_12078_ rbzero.color_sky\[1\] rbzero.color_floor\[1\] _04825_ vssd1 vssd1 vccd1 vccd1
+ _05267_ sky130_fd_sc_hd__mux2_1
XFILLER_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20285__152 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__inv_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15906_ _08555_ _08566_ _08564_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__a21o_1
X_11029_ rbzero.tex_b1\[22\] rbzero.tex_b1\[23\] _04303_ vssd1 vssd1 vccd1 vccd1 _04313_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16886_ _09906_ _09907_ vssd1 vssd1 vccd1 vccd1 _09908_ sky130_fd_sc_hd__nor2_1
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ _08919_ _08931_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__xor2_1
X_18625_ _02826_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__xnor2_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15768_ _08830_ _08861_ _08862_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18556_ rbzero.wall_tracer.rayAddendY\[-4\] _02527_ _02763_ _02766_ vssd1 vssd1 vccd1
+ vccd1 _00625_ sky130_fd_sc_hd__o22a_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17507_ _01797_ _01798_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__nor2_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14719_ _06575_ _07881_ _07888_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__o21a_1
X_18487_ _06092_ _06093_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__nor2_1
XFILLER_166_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15699_ _08787_ _08789_ _08792_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__and3_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17438_ _01727_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__and2_1
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _08148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _10311_ _10326_ vssd1 vssd1 vccd1 vccd1 _10387_ sky130_fd_sc_hd__or2_1
XFILLER_146_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20450__300 clknet_1_1__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__inv_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19108_ rbzero.spi_registers.texadd0\[8\] _03143_ vssd1 vssd1 vccd1 vccd1 _03153_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19039_ rbzero.map_overlay.i_othery\[2\] _03101_ vssd1 vssd1 vccd1 vccd1 _03112_
+ sky130_fd_sc_hd__or2_1
X_22050_ clknet_leaf_39_i_clk _01639_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21001_ clknet_leaf_100_i_clk _00590_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21903_ net429 _01492_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21834_ net360 _01423_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21765_ net291 _01354_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20716_ _03927_ _03924_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nor2_1
XFILLER_180_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21696_ net222 _01285_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20647_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__nand2_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ rbzero.tex_r1\[63\] net49 _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__mux2_1
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ _04534_ _04540_ _04543_ _03971_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a211o_1
XFILLER_178_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20578_ _09734_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13050_ _06120_ _06086_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or3_1
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12001_ _04826_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__buf_4
XFILLER_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ rbzero.wall_tracer.mapX\[6\] _09118_ vssd1 vssd1 vccd1 vccd1 _09778_ sky130_fd_sc_hd__xor2_1
XFILLER_98_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13952_ _06721_ _06708_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nand2_1
XFILLER_115_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ rbzero.map_rom.i_row\[4\] rbzero.wall_tracer.mapY\[5\] _06078_ vssd1 vssd1
+ vccd1 vccd1 _06079_ sky130_fd_sc_hd__o21a_1
X_16671_ _09749_ vssd1 vssd1 vccd1 vccd1 _09750_ sky130_fd_sc_hd__clkbuf_4
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13883_ _07011_ _07012_ _07014_ _07042_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and4_1
XFILLER_98_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15622_ _08715_ _08711_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__xor2_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18410_ _02637_ _02638_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__nand3_1
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12834_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__or2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19390_ _03116_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__buf_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _02574_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nand2_1
XFILLER_15_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15553_ _08634_ _08645_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__nor2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12765_ net38 net39 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__nor2_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14504_ _07045_ _07361_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__nor2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11716_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__buf_4
X_18272_ _02510_ _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__and2b_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15484_ _08383_ _08440_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__nor2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12696_ _05824_ _05829_ _05871_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a31o_2
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ _10021_ _10241_ vssd1 vssd1 vccd1 vccd1 _10243_ sky130_fd_sc_hd__or2_1
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14435_ _07586_ _07605_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__and2_1
X_11647_ _04835_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nand2_1
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput13 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_6
Xclkbuf_0__05700_ _05700_ vssd1 vssd1 vccd1 vccd1 clknet_0__05700_ sky130_fd_sc_hd__clkbuf_16
XFILLER_174_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17154_ _10171_ _10173_ vssd1 vssd1 vccd1 vccd1 _10174_ sky130_fd_sc_hd__nor2_1
XFILLER_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_190_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_4
XFILLER_167_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14366_ _07533_ _07535_ _07536_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__nand3_1
Xclkbuf_1_1__f__03792_ clknet_0__03792_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03792_
+ sky130_fd_sc_hd__clkbuf_16
X_11578_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand2_1
Xinput46 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_6
XFILLER_128_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16105_ _09197_ _09198_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__nand2_1
XFILLER_122_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13317_ _06413_ _06463_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__or2_1
X_17085_ _10076_ _10105_ vssd1 vssd1 vccd1 vccd1 _10106_ sky130_fd_sc_hd__xnor2_1
X_10529_ _04048_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14297_ _07357_ _07394_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__and2_1
XFILLER_182_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19675__55 clknet_1_1__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
X_16036_ _09077_ _09129_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13248_ rbzero.wall_tracer.visualWallDist\[8\] _04428_ _06324_ _06328_ vssd1 vssd1
+ vccd1 vccd1 _06419_ sky130_fd_sc_hd__o211a_1
XFILLER_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ _04443_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__nand2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_80_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _02196_ _02198_ _02194_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__o21a_1
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19726_ _03472_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
X_16938_ _09958_ _09959_ vssd1 vssd1 vccd1 vccd1 _09960_ sky130_fd_sc_hd__xor2_1
XFILLER_38_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _08616_ _09607_ _09890_ _09605_ vssd1 vssd1 vccd1 vccd1 _09891_ sky130_fd_sc_hd__a31o_1
XFILLER_168_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_95_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_203_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19588_ rbzero.spi_registers.new_texadd\[1\]\[11\] rbzero.spi_registers.spi_buffer\[11\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18539_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__nand2_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21550_ clknet_leaf_92_i_clk _01139_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20501_ clknet_1_0__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__buf_1
XFILLER_178_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21481_ net199 _01070_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22033_ clknet_leaf_67_i_clk _01622_ vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ rbzero.tex_g0\[30\] rbzero.tex_g0\[29\] _04226_ vssd1 vssd1 vccd1 vccd1 _04235_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20422__276 clknet_1_0__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__inv_2
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21817_ net343 _01406_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _05650_ _05704_ net12 _05730_ net11 vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__o2111a_1
X_21748_ net274 _01337_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11501_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__inv_2
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _05643_ _05658_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__nor2_1
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21679_ clknet_leaf_99_i_clk _01268_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ _07358_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ rbzero.spi_registers.texadd2\[3\] _04526_ rbzero.wall_hot\[0\] vssd1 vssd1
+ vccd1 vccd1 _04624_ sky130_fd_sc_hd__o21a_1
XFILLER_165_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _07206_ _07249_ _07205_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__or3b_1
XFILLER_165_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ _04454_ _04549_ _04552_ _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a31oi_1
XFILLER_4_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13102_ rbzero.wall_tracer.mapY\[8\] _06265_ _06266_ _06275_ vssd1 vssd1 vccd1 vccd1
+ _00388_ sky130_fd_sc_hd__a22o_1
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14082_ _06857_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__clkbuf_4
X_11294_ rbzero.spi_registers.texadd3\[8\] _04465_ _04455_ rbzero.spi_registers.texadd2\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__a22o_1
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17910_ _01818_ _01718_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__nor2_1
X_13033_ rbzero.wall_tracer.trackDistY\[4\] _06170_ rbzero.wall_tracer.trackDistY\[3\]
+ _06171_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__o221a_1
X_18890_ _03026_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17841_ _01997_ _01998_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__nand2_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17772_ _01940_ _01954_ _01952_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a21oi_1
X_14984_ _08101_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19511_ rbzero.spi_registers.got_new_texadd\[1\] _08117_ _03316_ _03383_ vssd1 vssd1
+ vccd1 vccd1 _00963_ sky130_fd_sc_hd__a31o_1
XFILLER_208_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13935_ _07104_ _07105_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__xor2_1
X_16723_ rbzero.wall_hot\[1\] rbzero.row_render.wall\[1\] _09760_ vssd1 vssd1 vccd1
+ vccd1 _09762_ sky130_fd_sc_hd__mux2_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19442_ rbzero.spi_registers.spi_buffer\[8\] rbzero.spi_registers.new_other\[8\]
+ _03338_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
X_16654_ _05069_ _09732_ vssd1 vssd1 vccd1 vccd1 _09737_ sky130_fd_sc_hd__and2_1
XFILLER_90_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13866_ _07018_ _07031_ _07036_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__o21ba_1
X_15605_ _08356_ _08697_ _08699_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__and3_1
XFILLER_179_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12817_ reg_gpout\[5\] clknet_1_0__leaf__05993_ net45 vssd1 vssd1 vccd1 vccd1 _05994_
+ sky130_fd_sc_hd__mux2_2
X_16585_ _09666_ _09674_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__xor2_1
X_19373_ rbzero.spi_registers.spi_done _02951_ _02929_ _02950_ vssd1 vssd1 vccd1 vccd1
+ _03306_ sky130_fd_sc_hd__and4b_1
XFILLER_37_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20397__253 clknet_1_0__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__inv_2
X_13797_ _06965_ _06964_ _06963_ _06957_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__a211oi_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15536_ _08599_ _08592_ _08598_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__a21oi_1
X_18324_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__or2_1
XFILLER_188_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12748_ _04643_ net28 _05922_ _05888_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a211oi_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18255_ _02502_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15467_ _08253_ _08276_ _08328_ _08327_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__or4_1
XFILLER_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ net44 _05845_ _05846_ _05848_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a311o_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17206_ _10087_ _10100_ _10225_ vssd1 vssd1 vccd1 vccd1 _10226_ sky130_fd_sc_hd__a21o_1
XFILLER_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14418_ _07582_ _07586_ _07587_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__nand3_1
XFILLER_198_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18186_ rbzero.wall_tracer.trackDistY\[7\] _02453_ _02336_ vssd1 vssd1 vccd1 vccd1
+ _02454_ sky130_fd_sc_hd__mux2_1
XFILLER_191_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15398_ _08483_ _08491_ _08492_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__a21o_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _10155_ _10156_ vssd1 vssd1 vccd1 vccd1 _10157_ sky130_fd_sc_hd__xor2_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14349_ _07481_ _07496_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17068_ _09974_ _09975_ _08431_ vssd1 vssd1 vccd1 vccd1 _10089_ sky130_fd_sc_hd__a21o_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16019_ _09108_ _09109_ _09112_ _09113_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__a31o_1
XFILLER_170_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20981_ clknet_leaf_64_i_clk _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21602_ clknet_leaf_91_i_clk _01191_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_181_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21533_ clknet_leaf_93_i_clk _01122_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21464_ net182 _01053_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21395_ clknet_leaf_4_i_clk _00984_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20346_ clknet_1_1__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__buf_1
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19654__36 clknet_1_0__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XFILLER_134_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22016_ clknet_leaf_69_i_clk _01605_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ rbzero.debug_overlay.playerY\[5\] _05101_ _05113_ rbzero.debug_overlay.playerY\[-4\]
+ _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a221o_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03795_ clknet_0__03795_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03795_
+ sky130_fd_sc_hd__clkbuf_16
X_13720_ _06682_ _06700_ _06784_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__and3_1
XFILLER_99_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10932_ _04262_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13651_ _06737_ _06725_ _06820_ _06821_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__nand4_1
X_10863_ _04214_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__clkbuf_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12602_ _05770_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__inv_2
XFILLER_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _09239_ _09337_ _09335_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__a21oi_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _06681_ _06725_ _06736_ _06739_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__a22o_1
X_10794_ rbzero.tex_g1\[6\] rbzero.tex_g1\[7\] _04188_ vssd1 vssd1 vccd1 vccd1 _04190_
+ sky130_fd_sc_hd__mux2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _08389_ _08415_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__or2b_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ _05711_ _05712_ _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__and3_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _02173_ _02259_ _02270_ _02326_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__o211a_1
XFILLER_185_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15252_ _08314_ _08346_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12464_ net4 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_80 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_80/HI o_rgb[5] sky130_fd_sc_hd__conb_1
XFILLER_32_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_91 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_91/HI o_rgb[20] sky130_fd_sc_hd__conb_1
X_14203_ _07371_ _07373_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__xnor2_1
X_11415_ rbzero.spi_registers.texadd2\[5\] _04537_ _04545_ rbzero.spi_registers.texadd1\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a22o_1
XFILLER_172_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ rbzero.debug_overlay.playerX\[-3\] _08254_ vssd1 vssd1 vccd1 vccd1 _08278_
+ sky130_fd_sc_hd__nand2_1
X_12395_ rbzero.tex_b1\[58\] _04914_ _04981_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a21o_1
XFILLER_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _06993_ _07303_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__or2_2
XFILLER_141_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11346_ rbzero.spi_registers.texadd3\[18\] _04526_ _04537_ rbzero.spi_registers.texadd2\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a22o_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19991_ rbzero.debug_overlay.playerY\[0\] _03617_ _03635_ _03630_ vssd1 vssd1 vccd1
+ vccd1 _01191_ sky130_fd_sc_hd__o211a_1
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _07218_ _07192_ _07235_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__a21oi_1
X_18942_ _02483_ _02481_ _03052_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
X_11277_ _04459_ rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__and2_1
XFILLER_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13016_ rbzero.wall_tracer.trackDistY\[-8\] _06186_ rbzero.wall_tracer.trackDistY\[-9\]
+ _06187_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o221a_1
X_18873_ _03017_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17824_ _02104_ _02112_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__xor2_1
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 rbzero.pov.spi_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17755_ _10288_ _09315_ _09195_ _01697_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__o22a_1
X_14967_ rbzero.wall_tracer.stepDistX\[-11\] _07867_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08093_ sky130_fd_sc_hd__mux2_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16706_ _09751_ vssd1 vssd1 vccd1 vccd1 _09757_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20405__260 clknet_1_0__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__inv_2
XFILLER_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13918_ _06726_ _06769_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__nor2_1
X_17686_ _10255_ _10256_ _10372_ _01975_ _01976_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__o41a_2
X_14898_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.trackDistX\[-9\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08044_ sky130_fd_sc_hd__mux2_1
XFILLER_165_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19425_ rbzero.spi_registers.got_new_leak _03118_ _03316_ _03336_ vssd1 vssd1 vccd1
+ vccd1 _00924_ sky130_fd_sc_hd__a31o_1
XFILLER_23_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _06772_ _06857_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__nor2_1
XFILLER_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16637_ _08148_ _09725_ _09726_ _04442_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__o211a_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ rbzero.spi_registers.new_floor\[5\] rbzero.spi_registers.got_new_floor _03097_
+ _04409_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a31o_1
X_16568_ _09656_ _09657_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__and2b_1
XFILLER_204_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18307_ rbzero.debug_overlay.vplaneX\[-7\] _02536_ vssd1 vssd1 vccd1 vccd1 _02545_
+ sky130_fd_sc_hd__nand2_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15519_ _08572_ _08613_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__xor2_1
X_16499_ _09463_ _09589_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__nand2_1
X_19287_ rbzero.spi_registers.texadd3\[11\] _03255_ vssd1 vssd1 vccd1 vccd1 _03257_
+ sky130_fd_sc_hd__or2_1
XFILLER_176_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18238_ _02493_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18169_ _02341_ _02437_ _02438_ _02339_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__o31a_1
XFILLER_190_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20200_ rbzero.spi_registers.new_texadd\[3\]\[15\] rbzero.spi_registers.spi_buffer\[15\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__mux2_1
XFILLER_85_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21180_ clknet_leaf_13_i_clk _00769_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20131_ _03722_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__and2b_1
Xclkbuf_0__03789_ _03789_ vssd1 vssd1 vccd1 vccd1 clknet_0__03789_ sky130_fd_sc_hd__clkbuf_16
X_20062_ rbzero.pov.ready_buffer\[29\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03683_
+ sky130_fd_sc_hd__and3_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ clknet_leaf_57_i_clk _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20895_ clknet_leaf_49_i_clk _00484_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21516_ clknet_leaf_82_i_clk _01105_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21447_ net165 _01036_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
X_20233__105 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__inv_2
XFILLER_163_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11200_ _04402_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12180_ _04941_ _05363_ _05367_ _04955_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a211o_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21378_ clknet_leaf_29_i_clk _00967_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11131_ _04366_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11062_ _04330_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15870_ _08912_ _08943_ _08964_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__a21oi_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _07866_ _07981_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__nand2_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _08889_ _08816_ _10093_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__or3_2
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _07822_ _07883_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__nand2_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _05148_ _05150_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or3_2
XFILLER_205_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03778_ clknet_0__03778_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03778_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _06866_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__xnor2_2
X_10915_ _04253_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] _10379_
+ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ _07850_ _07853_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__xnor2_1
X_11895_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__inv_2
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19210_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__clkbuf_4
XFILLER_204_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16422_ _09511_ _09512_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__nand2_1
X_13634_ _06790_ _06639_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__nor2_1
XFILLER_189_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ _04217_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16353_ _09442_ _09443_ _09415_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19141_ rbzero.spi_registers.new_texadd\[0\]\[22\] _03140_ _03171_ _03169_ vssd1
+ vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__o211a_1
XFILLER_73_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _06726_ _06727_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__or3b_2
XFILLER_34_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10777_ rbzero.tex_g1\[14\] rbzero.tex_g1\[15\] _04177_ vssd1 vssd1 vccd1 vccd1 _04181_
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15304_ _08392_ _08398_ _08158_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__mux2_4
XFILLER_9_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19072_ rbzero.spi_registers.new_mapd\[6\] _03120_ _03132_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00775_ sky130_fd_sc_hd__o211a_1
X_12516_ net9 _05697_ net5 _05640_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__and4b_1
X_16284_ _09271_ _09369_ _09375_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__a21o_1
XFILLER_160_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _06663_ _06599_ _06664_ _06665_ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__o32a_1
XFILLER_185_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ _08298_ _08327_ _08329_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__o21bai_1
X_18023_ _01818_ _10093_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor2_1
XFILLER_145_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ _05176_ _05550_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__and3b_4
XFILLER_154_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15166_ _08259_ _08260_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__nand2_1
XFILLER_114_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12378_ _04981_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__or2_1
XFILLER_158_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14117_ _07259_ _07275_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__a21oi_1
X_11329_ _04462_ _04517_ _04518_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__o211a_1
XFILLER_114_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19974_ rbzero.debug_overlay.playerY\[-5\] _03617_ _03623_ _03579_ vssd1 vssd1 vccd1
+ vccd1 _01186_ sky130_fd_sc_hd__o211a_1
X_15097_ rbzero.wall_tracer.visualWallDist\[-8\] _08160_ vssd1 vssd1 vccd1 vccd1 _08192_
+ sky130_fd_sc_hd__nor2_1
XFILLER_119_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18925_ _03044_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14048_ _06718_ _06727_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nor2_1
XFILLER_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18856_ _03008_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17807_ _02049_ _02057_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__nand2_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20329__191 clknet_1_1__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__inv_2
X_18787_ _02972_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15999_ _08367_ _08658_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__or2b_1
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _01995_ _02027_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17669_ _01804_ _01851_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a21oi_1
X_19408_ rbzero.spi_registers.got_new_floor _03118_ _03316_ _03326_ vssd1 vssd1 vccd1
+ vccd1 _00917_ sky130_fd_sc_hd__a31o_1
XFILLER_196_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20680_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03899_
+ sky130_fd_sc_hd__nand2_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19339_ rbzero.spi_registers.new_sky\[4\] rbzero.spi_registers.got_new_sky _03097_
+ _04409_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a31o_1
XFILLER_149_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21301_ clknet_leaf_29_i_clk _00890_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21232_ clknet_leaf_10_i_clk _00821_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21163_ clknet_leaf_95_i_clk _00752_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20114_ rbzero.pov.ready_buffer\[8\] _03663_ _03711_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01238_ sky130_fd_sc_hd__o211a_1
X_21094_ clknet_leaf_93_i_clk _00683_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20045_ net512 _03656_ _03673_ _03630_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__o211a_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21996_ net142 _01585_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ clknet_leaf_59_i_clk _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10700_ rbzero.tex_g1\[50\] rbzero.tex_g1\[51\] _04132_ vssd1 vssd1 vccd1 vccd1 _04140_
+ sky130_fd_sc_hd__mux2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ rbzero.row_render.size\[2\] _04446_ _04449_ rbzero.row_render.size\[1\] vssd1
+ vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__o22a_1
XFILLER_198_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20878_ clknet_leaf_36_i_clk _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ rbzero.tex_r0\[20\] rbzero.tex_r0\[19\] _04099_ vssd1 vssd1 vccd1 vccd1 _04104_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13350_ _06372_ _06503_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__xor2_4
X_10562_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _04066_ vssd1 vssd1 vccd1 vccd1 _04068_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ _05484_ _05485_ _05486_ _05190_ _04952_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__o221a_1
X_13281_ _06398_ _06400_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__and2_1
X_10493_ _04029_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__clkbuf_1
X_15020_ _08120_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
X_12232_ _04955_ _05405_ _05409_ _04887_ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a311o_1
XFILLER_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _04941_ _05350_ _04955_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__a21o_1
XFILLER_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11114_ _04357_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16971_ _09989_ _09991_ vssd1 vssd1 vccd1 vccd1 _09993_ sky130_fd_sc_hd__nand2_1
X_12094_ _03972_ _04418_ _04411_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__and3_1
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18710_ _02822_ _02794_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a21oi_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ _09014_ _09016_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__nor2_1
X_11045_ _04321_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ rbzero.debug_overlay.vplaneY\[-2\] _05129_ _02843_ vssd1 vssd1 vccd1 vccd1
+ _02845_ sky130_fd_sc_hd__o21ai_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _08944_ _08945_ _08947_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__a21o_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _07067_ _07855_ _07894_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__a21oi_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _02776_ _02777_ _02779_ _08134_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a31o_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _08873_ _08878_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__xor2_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ rbzero.wall_tracer.trackDistX\[2\] vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__inv_2
XFILLER_206_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17523_ _08814_ _09677_ _01814_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__or3_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ _05127_ _05105_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a21o_2
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _07827_ _07808_ _07818_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _10385_ _01746_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__xnor2_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _07836_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__inv_2
XFILLER_189_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ gpout0.hpos\[4\] _05061_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nor2_1
XFILLER_162_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16405_ _09378_ _09368_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__or2b_1
X_13617_ _06786_ _06787_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10829_ rbzero.tex_g0\[54\] rbzero.tex_g0\[53\] _04203_ vssd1 vssd1 vccd1 vccd1 _04208_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17385_ _08399_ _08618_ _01676_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__o21ai_1
X_14597_ _07718_ _07760_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__and2_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19124_ rbzero.spi_registers.new_texadd\[0\]\[14\] _03155_ _03162_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__o211a_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20517__361 clknet_1_1__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__inv_2
XFILLER_158_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16336_ rbzero.wall_tracer.visualWallDist\[-10\] _08149_ _09310_ vssd1 vssd1 vccd1
+ vccd1 _09428_ sky130_fd_sc_hd__and3_1
X_13548_ _06710_ _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__xor2_4
XFILLER_199_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16267_ _09260_ _09262_ _09358_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__o21ai_1
XFILLER_146_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19055_ rbzero.spi_registers.new_mapd\[10\] _03120_ _03123_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00767_ sky130_fd_sc_hd__o211a_1
XFILLER_199_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13479_ _06641_ _06644_ _06646_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__a211o_1
XFILLER_199_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _02285_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__xnor2_1
X_15218_ _06262_ _08308_ _08312_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__o21ai_4
XFILLER_173_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ _09038_ _09290_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__nand2_1
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _08242_ _08243_ _08157_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__mux2_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19957_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18908_ rbzero.pov.spi_buffer\[61\] rbzero.pov.ready_buffer\[61\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03036_ sky130_fd_sc_hd__mux2_1
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03457_ clknet_0__03457_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03457_
+ sky130_fd_sc_hd__clkbuf_16
X_19888_ rbzero.pov.ready _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and2_4
XFILLER_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18839_ _02999_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20262__131 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__inv_2
X_21850_ net376 _01439_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20801_ clknet_leaf_47_i_clk _00390_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21781_ net307 _01370_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20732_ _03936_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__buf_1
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20663_ _03882_ _03883_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__and3_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20594_ _03825_ _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nand2_1
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_104_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21215_ clknet_leaf_5_i_clk _00804_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21146_ clknet_leaf_99_i_clk _00735_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20345__206 clknet_1_0__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__inv_2
X_21077_ clknet_leaf_84_i_clk _00666_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20028_ _03654_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__clkbuf_4
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__nand2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04906_ _04988_ _04990_ _04920_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o211a_1
XFILLER_15_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ net34 vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ net505 _01568_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14520_ _07657_ _07656_ _07654_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__a21o_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _04827_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__buf_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _07599_ _07621_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__xor2_1
XFILLER_35_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11663_ _04835_ _04836_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or2_1
XFILLER_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _06566_ _06572_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and2_1
X_10614_ rbzero.tex_r0\[28\] rbzero.tex_r0\[27\] _04088_ vssd1 vssd1 vccd1 vccd1 _04095_
+ sky130_fd_sc_hd__mux2_1
X_17170_ _09670_ _09184_ _08813_ vssd1 vssd1 vccd1 vccd1 _10190_ sky130_fd_sc_hd__a21oi_2
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14382_ _07539_ _07548_ _07550_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__nor3_1
X_11594_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] _04783_ vssd1 vssd1 vccd1 vccd1
+ _04784_ sky130_fd_sc_hd__o21ai_2
XFILLER_70_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _09211_ _09213_ vssd1 vssd1 vccd1 vccd1 _09215_ sky130_fd_sc_hd__and2_1
XFILLER_70_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ _06372_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__xnor2_1
X_10545_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _04055_ vssd1 vssd1 vccd1 vccd1 _04059_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16052_ _08847_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13264_ _06425_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__nor2_1
X_10476_ _04020_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15003_ _08111_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
X_12215_ rbzero.tex_g1\[22\] _05236_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__or2_1
XFILLER_29_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13195_ _06299_ _06300_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__xor2_4
XFILLER_68_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19811_ rbzero.pov.spi_buffer\[43\] rbzero.pov.spi_buffer\[44\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03517_ sky130_fd_sc_hd__mux2_1
X_12146_ _05191_ _05331_ _05333_ _04953_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__o211a_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19742_ rbzero.pov.spi_buffer\[10\] rbzero.pov.spi_buffer\[11\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03481_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16954_ _09974_ _09975_ _08950_ vssd1 vssd1 vccd1 vccd1 _09976_ sky130_fd_sc_hd__a21o_1
X_12077_ _05017_ _05180_ _05265_ _04900_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__o211a_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11028_ _04312_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
X_15905_ _08659_ _08764_ _08997_ _08999_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__a22o_2
X_16885_ _09903_ _09905_ vssd1 vssd1 vccd1 vccd1 _09907_ sky130_fd_sc_hd__and2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18624_ _02827_ _02816_ _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__a21o_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _08920_ _08926_ _08930_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__o21a_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18555_ _02534_ _02764_ _02765_ _09745_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a31o_1
X_15767_ _08833_ _08860_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__nor2_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12979_ _04738_ _06088_ _06121_ rbzero.map_overlay.i_mapdy\[4\] _06154_ vssd1 vssd1
+ vccd1 vccd1 _06155_ sky130_fd_sc_hd__o221a_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17506_ _01794_ _01796_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__and2_1
XFILLER_205_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14718_ _06595_ _07887_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__or2_1
X_18486_ _06089_ _06265_ _02708_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a21oi_1
X_15698_ _08787_ _08789_ _08792_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__a21o_1
XFILLER_36_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _10096_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__xor2_1
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ _06613_ _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__or2_1
XANTENNA_16 _09747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_27 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 _05299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17368_ _10286_ _10303_ _10301_ vssd1 vssd1 vccd1 vccd1 _10386_ sky130_fd_sc_hd__a21o_1
XFILLER_186_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19107_ rbzero.spi_registers.new_texadd\[0\]\[7\] _03141_ _03152_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00790_ sky130_fd_sc_hd__o211a_1
X_16319_ _09293_ _09410_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__xnor2_1
X_17299_ _09528_ _09669_ vssd1 vssd1 vccd1 vccd1 _10318_ sky130_fd_sc_hd__nor2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19038_ rbzero.spi_registers.new_other\[1\] _03098_ _03109_ _03111_ vssd1 vssd1 vccd1
+ vccd1 _00762_ sky130_fd_sc_hd__o211a_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21000_ clknet_leaf_100_i_clk _00589_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21902_ net428 _01491_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21833_ net359 _01422_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21764_ net290 _01353_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20715_ _03927_ _03924_ _04442_ _04430_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__o211a_1
XFILLER_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21695_ net221 _01284_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20646_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03870_
+ sky130_fd_sc_hd__or2_1
XFILLER_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20577_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03813_
+ sky130_fd_sc_hd__or2_1
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12000_ rbzero.tex_r1\[10\] _05182_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__or2_1
XFILLER_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20269__137 clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__inv_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21129_ clknet_leaf_93_i_clk _00718_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13951_ _07120_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12902_ _06077_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__buf_2
XFILLER_189_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13882_ _07015_ _07041_ _07052_ _07014_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__o211a_1
X_16670_ _09748_ vssd1 vssd1 vccd1 vccd1 _09749_ sky130_fd_sc_hd__buf_4
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15621_ _08711_ _08715_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__or2b_1
X_12833_ _06005_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__nand2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__nand2_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _08301_ _08290_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__xnor2_1
X_12764_ net35 net34 vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nor2_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14503_ _07628_ _07670_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__xor2_1
X_15483_ _08502_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__xnor2_2
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18271_ _05111_ rbzero.wall_tracer.rayAddendX\[-5\] vssd1 vssd1 vccd1 vccd1 _02511_
+ sky130_fd_sc_hd__nand2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ clknet_1_0__leaf__04634_ _05845_ _05846_ _05873_ vssd1 vssd1 vccd1 vccd1
+ _05874_ sky130_fd_sc_hd__a31o_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _10021_ _10241_ vssd1 vssd1 vccd1 vccd1 _10242_ sky130_fd_sc_hd__nand2_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14434_ _07584_ _07585_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__or2_1
X_11646_ rbzero.row_render.size\[1\] rbzero.row_render.size\[0\] vssd1 vssd1 vccd1
+ vccd1 _04836_ sky130_fd_sc_hd__nor2_1
XFILLER_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_8
X_17153_ _10041_ _10048_ _10172_ vssd1 vssd1 vccd1 vccd1 _10173_ sky130_fd_sc_hd__a21oi_1
XFILLER_122_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14365_ _06942_ _07204_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__nor2_1
Xinput25 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_8
Xinput36 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_4
X_11577_ _04762_ _04766_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1__f__03791_ clknet_0__03791_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03791_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput47 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_4
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16104_ _08950_ _09186_ _09193_ _09196_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__o22ai_1
X_13316_ _06447_ _06436_ _06445_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__and3_1
XFILLER_196_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17084_ _10101_ _10104_ vssd1 vssd1 vccd1 vccd1 _10105_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10528_ rbzero.tex_r1\[2\] rbzero.tex_r1\[3\] _04046_ vssd1 vssd1 vccd1 vccd1 _04048_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14296_ _07413_ _07466_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__nor2_1
XFILLER_183_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16035_ _08335_ _08618_ vssd1 vssd1 vccd1 vccd1 _09129_ sky130_fd_sc_hd__nor2_1
XFILLER_182_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _06393_ _06406_ _06408_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__nand3_1
X_10459_ _04011_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13178_ _06346_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12129_ _04923_ _05313_ _05316_ _04953_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__o211a_1
X_17986_ _02221_ _02222_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__o22a_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20480__327 clknet_1_1__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__inv_2
XFILLER_46_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19725_ rbzero.pov.spi_buffer\[2\] rbzero.pov.spi_buffer\[3\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
X_16937_ _09044_ _09046_ _09406_ vssd1 vssd1 vccd1 vccd1 _09959_ sky130_fd_sc_hd__a21o_1
XFILLER_133_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16868_ _09687_ vssd1 vssd1 vccd1 vccd1 _09890_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18607_ _02796_ _02811_ _02810_ _02809_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__o211ai_2
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _08228_ _08696_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__or3b_1
XFILLER_203_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19587_ _03422_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__clkbuf_1
X_16799_ _09825_ _09826_ _09827_ vssd1 vssd1 vccd1 vccd1 _09829_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18538_ _02747_ _02748_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__o21ba_1
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18469_ _02694_ _02681_ _02685_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a21oi_1
X_20374__232 clknet_1_0__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__inv_2
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21480_ net198 _01069_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22032_ clknet_leaf_54_i_clk _01621_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21816_ net342 _01405_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21747_ net273 _01336_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _04684_ _04685_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__and3_1
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12480_ _05661_ _05640_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nand2_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21678_ clknet_leaf_1_i_clk _01267_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ rbzero.spi_registers.texadd3\[3\] _04457_ _04545_ rbzero.spi_registers.texadd1\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a22o_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20629_ _03849_ _03852_ _03850_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__o21ai_1
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ _06775_ _07310_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__nand2_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _04454_ _04552_ _04553_ _04549_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a22oi_1
XFILLER_192_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13101_ _06272_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__xor2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_i_clk clknet_1_0_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14081_ _06942_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__clkbuf_4
X_11293_ rbzero.texu_hot\[3\] _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__nand2_1
X_13032_ rbzero.wall_tracer.trackDistY\[3\] _06171_ rbzero.wall_tracer.trackDistY\[2\]
+ _06172_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__a221o_1
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17840_ _02127_ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__xor2_1
XFILLER_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17771_ _02041_ _02060_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14983_ rbzero.wall_tracer.stepDistX\[-3\] _07971_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08101_ sky130_fd_sc_hd__mux2_1
XFILLER_87_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19510_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__buf_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16722_ _09761_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__clkbuf_1
X_13934_ _06971_ _06930_ _06928_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__o21ba_1
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19441_ _03345_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16653_ _05075_ _09730_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__nor2_1
X_13865_ _07034_ _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__nor2_1
X_15604_ _08359_ _08698_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ _05632_ _05940_ _05943_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__o31a_2
X_19372_ rbzero.spi_registers.new_vshift\[5\] _03297_ _03305_ _03302_ vssd1 vssd1
+ vccd1 vccd1 _00902_ sky130_fd_sc_hd__o211a_1
XFILLER_76_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16584_ _09663_ _09673_ vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__xor2_1
X_13796_ _06960_ _06961_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__or2_1
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18323_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__nand2_1
XFILLER_72_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15535_ _08599_ _08592_ _08598_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__and3_1
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ net55 _05910_ _05920_ net53 _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a221o_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ rbzero.spi_registers.new_texadd\[2\]\[16\] rbzero.spi_registers.spi_buffer\[16\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_187_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15466_ _08559_ _08560_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__xnor2_1
X_12678_ net25 _05835_ _05850_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a31o_1
XFILLER_187_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17205_ _10097_ _10099_ vssd1 vssd1 vccd1 vccd1 _10225_ sky130_fd_sc_hd__nor2_1
X_11629_ _04812_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__or2_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14417_ _07582_ _07586_ _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__a21o_1
X_18185_ _02451_ _02452_ _02083_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__o21ai_1
X_15397_ _08486_ _08490_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__nor2_1
XFILLER_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17136_ _08952_ _09491_ _10030_ _10032_ vssd1 vssd1 vccd1 vccd1 _10156_ sky130_fd_sc_hd__o31a_1
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14348_ _07475_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17067_ _09167_ _09560_ vssd1 vssd1 vccd1 vccd1 _10088_ sky130_fd_sc_hd__or2_1
X_14279_ _07448_ _07449_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__or2_1
XFILLER_83_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16018_ _09110_ _09111_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__and2_1
XFILLER_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _02184_ _02185_ _02254_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__and3_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_100_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20980_ clknet_leaf_64_i_clk _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19639_ rbzero.pov.spi_counter\[5\] _03451_ _03440_ vssd1 vssd1 vccd1 vccd1 _03455_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21601_ clknet_leaf_91_i_clk _01190_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21532_ clknet_leaf_93_i_clk _01121_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21463_ net181 _01052_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21394_ clknet_leaf_2_i_clk _00983_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22015_ clknet_leaf_48_i_clk _01604_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _04656_ gpout0.vpos\[4\] gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _05169_
+ sky130_fd_sc_hd__or3b_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03794_ clknet_0__03794_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03794_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ rbzero.tex_g0\[6\] rbzero.tex_g0\[5\] _04259_ vssd1 vssd1 vccd1 vccd1 _04262_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ _04225_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
X_13650_ _06728_ _06738_ _06759_ _06700_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a22o_1
XFILLER_204_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _04687_ _05644_ _05645_ _04642_ _05763_ _05770_ vssd1 vssd1 vccd1 vccd1 _05781_
+ sky130_fd_sc_hd__mux4_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13581_ _06707_ _06741_ _06744_ _06746_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a32o_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _04189_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__clkbuf_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15320_ _08411_ _08412_ _08413_ _08414_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12532_ net14 net15 vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nor2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15251_ _08325_ _08337_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__nor2_1
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12463_ _04648_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__buf_2
XFILLER_173_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_81 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_81/HI o_rgb[8] sky130_fd_sc_hd__conb_1
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14202_ _07318_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__nand2_1
X_11414_ _03970_ _04603_ _04604_ _04605_ _04575_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
Xtop_ew_algofoogle_92 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_92/HI o_rgb[21] sky130_fd_sc_hd__conb_1
XFILLER_32_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15182_ rbzero.debug_overlay.playerX\[-3\] _08254_ vssd1 vssd1 vccd1 vccd1 _08277_
+ sky130_fd_sc_hd__or2_1
X_12394_ rbzero.tex_b1\[59\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__and3_1
XFILLER_158_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14133_ _07252_ _07253_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__or3_1
X_20511__356 clknet_1_1__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__inv_2
X_11345_ _04456_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__clkbuf_4
X_19990_ rbzero.pov.ready_buffer\[53\] _03570_ _03610_ _03634_ vssd1 vssd1 vccd1 vccd1
+ _03635_ sky130_fd_sc_hd__a211o_1
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_94_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _07233_ _07234_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__nand2_1
X_18941_ _03054_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
X_11276_ rbzero.spi_registers.texadd1\[12\] _04461_ vssd1 vssd1 vccd1 vccd1 _04468_
+ sky130_fd_sc_hd__and2_1
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13015_ rbzero.wall_tracer.trackDistY\[-9\] _06187_ rbzero.wall_tracer.trackDistY\[-10\]
+ _06188_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__a221o_1
X_18872_ rbzero.pov.spi_buffer\[44\] rbzero.pov.ready_buffer\[44\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17823_ _02110_ _02111_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__nor2_1
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 rbzero.pov.ready_buffer\[43\] vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17754_ _10288_ _09195_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__nor2_1
X_14966_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__buf_4
XFILLER_48_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ rbzero.traced_texa\[-1\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__a22o_1
X_13917_ _06866_ _06873_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a21oi_1
X_17685_ _01975_ _01755_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__or2b_1
X_14897_ _08036_ _08041_ _08043_ _01633_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__o211a_1
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19424_ _03329_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__inv_2
X_16636_ rbzero.texu_hot\[5\] _08145_ vssd1 vssd1 vccd1 vccd1 _09726_ sky130_fd_sc_hd__or2_1
X_13848_ _06754_ _06726_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__nor2_1
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19355_ rbzero.spi_registers.new_floor\[4\] _03289_ _03295_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00895_ sky130_fd_sc_hd__o211a_1
X_16567_ _09654_ _09655_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__nand2_1
XFILLER_210_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__05993_ clknet_0__05993_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05993_
+ sky130_fd_sc_hd__clkbuf_16
X_13779_ _06903_ _06948_ _06742_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__a21bo_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18306_ rbzero.debug_overlay.vplaneX\[-7\] _02536_ vssd1 vssd1 vccd1 vccd1 _02544_
+ sky130_fd_sc_hd__or2_1
X_15518_ _08603_ _08612_ _08601_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19286_ rbzero.spi_registers.new_texadd\[3\]\[10\] _03254_ _03256_ _03252_ vssd1
+ vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__o211a_1
X_16498_ _09587_ _09588_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__and2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18237_ rbzero.spi_registers.new_texadd\[2\]\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _02479_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_198_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15449_ _08534_ _08536_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__xor2_1
XFILLER_157_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18168_ _02434_ _02435_ _02436_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__o21a_1
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _10137_ _10131_ _10135_ _10136_ vssd1 vssd1 vccd1 vccd1 _10139_ sky130_fd_sc_hd__o211ai_2
XFILLER_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18099_ rbzero.wall_tracer.trackDistY\[-5\] _02378_ _02339_ vssd1 vssd1 vccd1 vccd1
+ _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_144_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20130_ _03973_ _09727_ _03721_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a31o_1
X_20486__333 clknet_1_0__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__inv_2
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03788_ _03788_ vssd1 vssd1 vccd1 vccd1 clknet_0__03788_ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20061_ rbzero.pov.ready_buffer\[28\] _03656_ _03682_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01214_ sky130_fd_sc_hd__o211a_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ clknet_leaf_57_i_clk _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ clknet_leaf_49_i_clk _00483_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21515_ clknet_leaf_81_i_clk _01104_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21446_ net164 _01035_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21377_ clknet_leaf_29_i_clk _00966_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _04362_ vssd1 vssd1 vccd1 vccd1 _04366_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ rbzero.tex_b1\[7\] rbzero.tex_b1\[8\] _04325_ vssd1 vssd1 vccd1 vccd1 _04330_
+ sky130_fd_sc_hd__mux2_1
XFILLER_192_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _06602_ _07897_ _07980_ _06655_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__a22oi_4
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _07913_ _07916_ _07918_ _06470_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__a211o_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ rbzero.debug_overlay.facingX\[10\] _05105_ _05115_ rbzero.debug_overlay.facingX\[0\]
+ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a221o_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03777_ clknet_0__03777_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03777_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06867_ _06872_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ rbzero.tex_g0\[14\] rbzero.tex_g0\[13\] _04248_ vssd1 vssd1 vccd1 vccd1 _04253_
+ sky130_fd_sc_hd__mux2_1
X_17470_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__and2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ _05061_ _05077_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or2_1
X_14682_ _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__inv_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16421_ _09485_ _09486_ _09510_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__nand3_1
X_10845_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _04215_ vssd1 vssd1 vccd1 vccd1 _04217_
+ sky130_fd_sc_hd__mux2_1
X_13633_ _06789_ _06794_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__xor2_1
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19140_ rbzero.spi_registers.texadd0\[22\] _03142_ vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__or2_1
X_16352_ _09415_ _09442_ _09443_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__and3_1
X_10776_ _04180_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13564_ _06728_ _06708_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__and3_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _08144_ _08394_ _08397_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__o21ai_2
XFILLER_201_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19071_ rbzero.map_overlay.i_mapdy\[2\] _03122_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__or2_1
X_12515_ _05693_ _05694_ _05695_ _05696_ net8 vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a32o_1
X_16283_ _09373_ _09374_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__nand2_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13495_ _06498_ _06582_ _06603_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__mux2_1
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ _02237_ _02302_ _02307_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a31o_1
XFILLER_201_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ _08276_ _08328_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__nor2_1
X_12446_ _05047_ _04744_ _05547_ _05630_ _04650_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a311o_1
XFILLER_173_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12377_ rbzero.tex_b1\[47\] rbzero.tex_b1\[46\] _04893_ vssd1 vssd1 vccd1 vccd1 _05562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15165_ rbzero.debug_overlay.playerY\[-5\] _08221_ rbzero.debug_overlay.playerY\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _04519_ _04461_ _04458_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21oi_1
X_14116_ _07276_ _07278_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__and2b_1
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19973_ rbzero.pov.ready_buffer\[48\] _03438_ _03610_ _03622_ vssd1 vssd1 vccd1 vccd1
+ _03623_ sky130_fd_sc_hd__a211o_1
X_15096_ _08189_ _08190_ _06075_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__mux2_1
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ rbzero.pov.spi_buffer\[69\] rbzero.pov.ready_buffer\[69\] _02967_ vssd1 vssd1
+ vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XFILLER_171_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14047_ _07127_ _07180_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__or2b_1
X_11259_ _04446_ _04447_ _04448_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a31o_1
XFILLER_141_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18855_ rbzero.pov.spi_buffer\[36\] rbzero.pov.ready_buffer\[36\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17806_ _02091_ _02094_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__xor2_1
XFILLER_83_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18786_ rbzero.pov.spi_buffer\[3\] rbzero.pov.ready_buffer\[3\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02972_ sky130_fd_sc_hd__mux2_1
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15998_ _08625_ _09092_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17737_ _02025_ _02026_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__nand2_1
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14949_ _08065_ _08079_ _08080_ _08061_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__o211a_1
XFILLER_209_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _01848_ _01850_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__nor2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19407_ _03319_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__inv_2
X_16619_ _09705_ _09707_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__nand2_1
X_17599_ _09520_ _09621_ _01775_ _01777_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__o31a_1
XFILLER_126_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19338_ rbzero.spi_registers.new_sky\[3\] _03280_ _03285_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00888_ sky130_fd_sc_hd__o211a_1
XFILLER_176_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19269_ rbzero.spi_registers.new_texadd\[3\]\[3\] _03240_ _03246_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00858_ sky130_fd_sc_hd__o211a_1
XFILLER_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21300_ clknet_leaf_31_i_clk _00889_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_129_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21231_ clknet_leaf_12_i_clk _00820_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21162_ clknet_leaf_94_i_clk _00751_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20113_ rbzero.debug_overlay.vplaneY\[-1\] _03685_ vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__or2_1
X_21093_ clknet_leaf_93_i_clk _00682_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20044_ rbzero.debug_overlay.facingX\[10\] _03658_ vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__or2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_0_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ net141 _01584_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20540__382 clknet_1_1__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__inv_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ clknet_leaf_59_i_clk _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ clknet_leaf_20_i_clk _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10630_ _04103_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ _04067_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12300_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _05009_ vssd1 vssd1 vccd1 vccd1 _05486_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13280_ _06449_ _06450_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__xnor2_1
X_10492_ rbzero.tex_r1\[19\] rbzero.tex_r1\[20\] _04024_ vssd1 vssd1 vccd1 vccd1 _04029_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _05411_ _05413_ _05415_ _05417_ _04902_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__o221a_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21429_ clknet_leaf_96_i_clk _01018_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ _05348_ _05349_ _05191_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__mux2_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11113_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _04351_ vssd1 vssd1 vccd1 vccd1 _04357_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16970_ _09989_ _09991_ vssd1 vssd1 vccd1 vccd1 _09992_ sky130_fd_sc_hd__or2_1
X_12093_ _04657_ _04589_ _05280_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a31o_1
XFILLER_7_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15921_ _08276_ _08535_ _08558_ _09015_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__o31a_1
X_11044_ rbzero.tex_b1\[15\] rbzero.tex_b1\[16\] _04314_ vssd1 vssd1 vccd1 vccd1 _04321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ rbzero.debug_overlay.vplaneY\[-2\] _05129_ _02843_ vssd1 vssd1 vccd1 vccd1
+ _02844_ sky130_fd_sc_hd__or3_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _08696_ _08733_ _08946_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__and3b_1
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14803_ _07894_ _07926_ _07927_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__a21o_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _02776_ _02777_ _02779_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _08874_ _08877_ _08875_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__a21oi_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ rbzero.wall_tracer.trackDistX\[3\] vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__inv_2
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _09528_ _09559_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__or2_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14734_ _06619_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__buf_2
XFILLER_205_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ rbzero.debug_overlay.vplaneY\[-3\] _05110_ _05128_ _05131_ _05134_ vssd1
+ vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__a2111o_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__and2b_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _07834_ _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__and2_1
XFILLER_205_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _04640_ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__or2_1
X_16404_ _09487_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__xnor2_1
X_13616_ _06772_ _06729_ _06717_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__mux2_1
X_10828_ _04207_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__clkbuf_1
X_17384_ _08399_ _08618_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or3_1
X_20551__12 clknet_1_0__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
XFILLER_125_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14596_ _07763_ _07766_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__nand2_1
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19123_ rbzero.spi_registers.texadd0\[14\] _03156_ vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__or2_1
XFILLER_201_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16335_ _08471_ _09311_ _09426_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__nand3_1
Xclkbuf_1_1__f__05761_ clknet_0__05761_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05761_
+ sky130_fd_sc_hd__clkbuf_16
X_13547_ _06717_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10759_ _04171_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19054_ rbzero.map_overlay.i_mapdx\[0\] _03122_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__or2_1
X_16266_ _09244_ _09263_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__nand2_1
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _06537_ _06539_ _06647_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__a22o_1
XFILLER_173_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18005_ _02289_ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15217_ _08310_ _08311_ _08158_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__mux2_1
X_12429_ rbzero.tex_b1\[26\] _04908_ _04817_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a21o_1
XFILLER_127_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16197_ _09043_ _09046_ _08910_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__a21oi_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15148_ rbzero.wall_tracer.visualWallDist\[-5\] _08160_ vssd1 vssd1 vccd1 vccd1 _08243_
+ sky130_fd_sc_hd__or2_1
XFILLER_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19956_ net41 _03557_ _03095_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o21ai_4
X_15079_ rbzero.side_hot _06353_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__nand2_1
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18907_ _03035_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19887_ net41 net40 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__nor2_1
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18838_ rbzero.pov.spi_buffer\[28\] rbzero.pov.ready_buffer\[28\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18769_ _02952_ _02959_ _02960_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__nor3_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20800_ clknet_leaf_47_i_clk _00389_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21780_ net306 _01369_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20731_ _03728_ clknet_1_1__leaf__05993_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__and2_2
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20662_ _03877_ _03881_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nand2_1
XFILLER_196_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20593_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03826_
+ sky130_fd_sc_hd__nand2_1
XFILLER_104_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21214_ clknet_leaf_5_i_clk _00803_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21145_ clknet_leaf_1_i_clk _00734_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_160_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21076_ clknet_leaf_82_i_clk _00665_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20027_ rbzero.pov.ready_buffer\[36\] _03656_ _03662_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01200_ sky130_fd_sc_hd__o211a_1
XFILLER_150_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _04947_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _05952_ _05949_ _05955_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__o211a_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ net504 _01567_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _04906_ _04911_ _04916_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__o211a_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20929_ clknet_leaf_54_i_clk _00518_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _07601_ _07619_ _07620_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__a21oi_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _04838_ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
XFILLER_23_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ _06569_ _06538_ _06570_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a22o_1
X_10613_ _04094_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11593_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] rbzero.texV\[1\] rbzero.traced_texVinit\[1\]
+ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a221o_1
XFILLER_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14381_ _07498_ _07517_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__xnor2_1
X_16120_ _09211_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__nor2_1
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10544_ _04058_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13332_ _06370_ _06415_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__nand2_2
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16051_ _09031_ _09026_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__or2b_1
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10475_ rbzero.tex_r1\[27\] rbzero.tex_r1\[28\] _04013_ vssd1 vssd1 vccd1 vccd1 _04020_
+ sky130_fd_sc_hd__mux2_1
X_13263_ _06433_ rbzero.wall_tracer.visualWallDist\[9\] _04428_ _04444_ vssd1 vssd1
+ vccd1 vccd1 _06434_ sky130_fd_sc_hd__or4_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15002_ rbzero.wall_tracer.stepDistX\[6\] _08018_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08111_ sky130_fd_sc_hd__mux2_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12214_ _04903_ _05387_ _05391_ _04958_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a311o_1
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ rbzero.wall_tracer.rcp_sel\[0\] _06362_ _06363_ _06364_ vssd1 vssd1 vccd1
+ vccd1 _06365_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_194_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _05199_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__or2_1
X_19810_ _03516_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ _04810_ _05207_ _05225_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a31o_1
X_16953_ rbzero.wall_tracer.stepDistX\[9\] _09045_ vssd1 vssd1 vccd1 vccd1 _09975_
+ sky130_fd_sc_hd__nand2_2
X_19741_ _03480_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11027_ rbzero.tex_b1\[23\] rbzero.tex_b1\[24\] _04303_ vssd1 vssd1 vccd1 vccd1 _04312_
+ sky130_fd_sc_hd__mux2_1
X_15904_ _08659_ _08998_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__xnor2_2
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16884_ _09903_ _09905_ vssd1 vssd1 vccd1 vccd1 _09906_ sky130_fd_sc_hd__nor2_1
XFILLER_65_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18623_ _02818_ _02817_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__and2b_1
XFILLER_77_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _08928_ _08929_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__nand2_1
XFILLER_65_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18554_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__nand2_1
XFILLER_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15766_ _08833_ _08860_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__xor2_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ rbzero.map_overlay.i_mapdy\[3\] rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1
+ _06154_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _01794_ _01796_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__nor2_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14717_ _07883_ _07886_ _06584_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__mux2_1
X_18485_ _06111_ _08124_ _02704_ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__o211a_1
X_11929_ _05085_ _05116_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__nor2_4
X_15697_ _08529_ _08733_ _08790_ _08791_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__a31o_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17436_ _09167_ _01728_ _10342_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__mux2_2
X_14648_ _07790_ _07792_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _09747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17367_ _10383_ _10384_ vssd1 vssd1 vccd1 vccd1 _10385_ sky130_fd_sc_hd__nor2_1
X_14579_ _07423_ _07361_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__nor2_1
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19106_ rbzero.spi_registers.texadd0\[7\] _03143_ vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__or2_1
X_16318_ _08369_ _09037_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__nor2_1
XFILLER_158_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20292__158 clknet_1_0__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__inv_2
X_17298_ _10314_ _10316_ vssd1 vssd1 vccd1 vccd1 _10317_ sky130_fd_sc_hd__and2_1
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19037_ _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__buf_2
X_16249_ _09222_ _09224_ _09340_ _09341_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__or4bb_1
XFILLER_174_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19939_ rbzero.pov.ready_buffer\[70\] _03438_ _03558_ _03596_ vssd1 vssd1 vccd1 vccd1
+ _03597_ sky130_fd_sc_hd__a211o_1
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21901_ net427 _01490_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21832_ net358 _01421_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21763_ net289 _01352_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
X_20714_ _04436_ _04437_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__nand2_1
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21694_ net220 _01283_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20645_ _03734_ _03868_ _03869_ _03740_ rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1
+ _01611_ sky130_fd_sc_hd__a32o_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03812_
+ sky130_fd_sc_hd__nand2_1
X_20351__211 clknet_1_0__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__inv_2
XFILLER_20_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21128_ clknet_leaf_93_i_clk _00717_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21059_ clknet_leaf_98_i_clk _00648_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13950_ _06707_ _07078_ _06759_ _06722_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o22a_1
XFILLER_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12901_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13881_ _07038_ _07039_ _07048_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a211oi_1
XFILLER_189_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15620_ _08672_ _08712_ _08713_ _08714_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12832_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__nor2_1
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _08634_ _08645_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__xor2_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ net37 net36 vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__or2_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _07671_ _07672_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__and2_1
X_11714_ _04891_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__buf_4
X_18270_ _05111_ rbzero.wall_tracer.rayAddendX\[-5\] vssd1 vssd1 vccd1 vccd1 _02510_
+ sky130_fd_sc_hd__nor2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _08404_ _08457_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__nor2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ gpout3.clk_div\[1\] _05846_ _05847_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_
+ sky130_fd_sc_hd__a31o_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17221_ _10239_ _10240_ vssd1 vssd1 vccd1 vccd1 _10241_ sky130_fd_sc_hd__xor2_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14433_ _07558_ _07563_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11645_ rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__inv_2
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03459_ clknet_0__03459_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03459_
+ sky130_fd_sc_hd__clkbuf_16
X_17152_ _09936_ _09938_ _10047_ vssd1 vssd1 vccd1 vccd1 _10172_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14364_ _06741_ _07310_ _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__a21o_1
Xinput15 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__03790_ clknet_0__03790_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03790_
+ sky130_fd_sc_hd__clkbuf_16
X_11576_ rbzero.texV\[5\] _04765_ _04763_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a21oi_2
Xinput26 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_4
XFILLER_183_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16103_ _08441_ _09186_ _09193_ _09196_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__or4_1
XFILLER_155_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput48 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_8
X_13315_ _06453_ _06460_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__xnor2_4
X_10527_ _04047_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__clkbuf_1
X_17083_ _10102_ _10103_ _09983_ _09984_ _09964_ vssd1 vssd1 vccd1 vccd1 _10104_ sky130_fd_sc_hd__a32o_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14295_ _07414_ _07461_ _07465_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__o21a_1
XFILLER_202_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _09008_ _08553_ _09007_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__or3_1
X_10458_ rbzero.tex_r1\[35\] rbzero.tex_r1\[36\] _04002_ vssd1 vssd1 vccd1 vccd1 _04011_
+ sky130_fd_sc_hd__mux2_1
X_13246_ _06336_ _06338_ _06344_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__a21o_1
XFILLER_170_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ _06288_ _06347_ _06311_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__a21oi_1
X_10389_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12128_ _04982_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__or2_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17985_ _02251_ _02252_ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16936_ _09667_ _09957_ vssd1 vssd1 vccd1 vccd1 _09958_ sky130_fd_sc_hd__xnor2_1
X_12059_ rbzero.tex_r1\[60\] _04935_ _05195_ _05246_ _05247_ vssd1 vssd1 vccd1 vccd1
+ _05248_ sky130_fd_sc_hd__a311o_1
X_19724_ _03471_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19655_ clknet_1_0__leaf__03457_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__buf_1
X_16867_ _09889_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15818_ _08911_ _08912_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__xnor2_1
X_18606_ _02809_ _02810_ _02811_ _02796_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a211o_1
X_19586_ rbzero.spi_registers.new_texadd\[1\]\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__mux2_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16798_ _09825_ _09826_ _09827_ vssd1 vssd1 vccd1 vccd1 _09828_ sky130_fd_sc_hd__and3_1
XFILLER_19_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18537_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__and2_1
X_15749_ _08734_ _08233_ _08472_ _08457_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__or4_1
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ _02598_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__inv_2
XFILLER_179_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17419_ _01704_ _01710_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__or2_1
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18399_ _02616_ _02621_ _02628_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__or3_1
XFILLER_187_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22031_ clknet_leaf_41_i_clk _01620_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21815_ net341 _01404_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21746_ net272 _01335_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21677_ clknet_leaf_99_i_clk _01266_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ rbzero.spi_registers.texadd0\[2\] _04535_ _04621_ _03969_ vssd1 vssd1 vccd1
+ vccd1 _04622_ sky130_fd_sc_hd__o211a_1
XFILLER_165_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20628_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03855_
+ sky130_fd_sc_hd__nand2_1
XFILLER_177_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11361_ _04454_ _04544_ _04548_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or3_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13100_ _06100_ _06099_ _06267_ _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a31o_1
XFILLER_192_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ _07206_ _07249_ _07205_ _07250_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__o31a_1
X_11292_ rbzero.spi_registers.texadd0\[9\] _04467_ _04482_ _04483_ vssd1 vssd1 vccd1
+ vccd1 _04484_ sky130_fd_sc_hd__o22a_1
XFILLER_106_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _06178_ _06181_ _06196_ _06201_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__o41a_1
XFILLER_65_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17770_ _02042_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14982_ _08100_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16721_ rbzero.wall_hot\[0\] rbzero.row_render.wall\[0\] _09760_ vssd1 vssd1 vccd1
+ vccd1 _09761_ sky130_fd_sc_hd__mux2_1
X_13933_ _07101_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19440_ rbzero.spi_registers.spi_buffer\[7\] rbzero.spi_registers.new_other\[7\]
+ _03338_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__mux2_1
XFILLER_75_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16652_ _09736_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__clkbuf_1
X_13864_ _07018_ _07031_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15603_ _08346_ _08356_ _08360_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__a21oi_1
X_12815_ net39 _05961_ _05975_ _05981_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a311o_2
X_19371_ rbzero.spi_registers.vshift\[5\] _03298_ vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__or2_1
X_16583_ _09557_ _09667_ _09672_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__a21oi_1
X_13795_ _06957_ _06963_ _06964_ _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o211a_2
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18322_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__or2_1
XFILLER_16_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15534_ _08603_ _08612_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__xnor2_1
X_20358__217 clknet_1_0__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__inv_2
XFILLER_128_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ net52 _05921_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__and2_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18253_ _02501_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__clkbuf_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _08276_ _08340_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__or2_1
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12677_ _05824_ _05829_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a31o_1
XFILLER_169_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17204_ _10213_ _10223_ vssd1 vssd1 vccd1 vccd1 _10224_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ _07544_ _07546_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ _04814_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nand2_1
X_18184_ _02449_ _02450_ _09866_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a21o_1
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15396_ _08486_ _08490_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__xor2_2
XFILLER_156_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17135_ _10153_ _10154_ vssd1 vssd1 vccd1 vccd1 _10155_ sky130_fd_sc_hd__nand2_1
XFILLER_184_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ _07498_ _07517_ _07515_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _04749_ sky130_fd_sc_hd__nand2_1
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17066_ _10078_ _10086_ vssd1 vssd1 vccd1 vccd1 _10087_ sky130_fd_sc_hd__xor2_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14278_ _07206_ _07361_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__nor2_1
XFILLER_48_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _09110_ _09111_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__or2_1
X_13229_ _04428_ _06044_ _06045_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a31o_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17968_ _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__inv_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16919_ _08813_ _09176_ vssd1 vssd1 vccd1 vccd1 _09941_ sky130_fd_sc_hd__nor2_1
X_17899_ _02104_ _02112_ _02110_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a21o_1
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19638_ rbzero.pov.spi_counter\[5\] _03451_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and2_1
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19569_ rbzero.spi_registers.new_texadd\[1\]\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21600_ clknet_leaf_91_i_clk _01189_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_209_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20298__164 clknet_1_1__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__inv_2
XFILLER_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21531_ clknet_leaf_97_i_clk _01120_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21462_ net180 _01051_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21393_ clknet_leaf_2_i_clk _00982_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22014_ clknet_leaf_69_i_clk _01603_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20463__312 clknet_1_0__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__inv_2
XFILLER_76_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03793_ clknet_0__03793_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03793_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ _04261_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10861_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _04215_ vssd1 vssd1 vccd1 vccd1 _04225_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ net17 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__inv_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ _06687_ _06750_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__nor2_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ rbzero.tex_g1\[7\] rbzero.tex_g1\[8\] _04188_ vssd1 vssd1 vccd1 vccd1 _04189_
+ sky130_fd_sc_hd__mux2_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12531_ net11 _05704_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__and2_1
X_21729_ net255 _01318_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _08340_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__nor2_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _04653_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__buf_2
XFILLER_40_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14201_ _07316_ _07249_ _07317_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__o21bai_1
Xtop_ew_algofoogle_82 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_82/HI o_rgb[9] sky130_fd_sc_hd__conb_1
X_11413_ _03970_ _04498_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__nor2_1
Xtop_ew_algofoogle_93 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_93/HI zeros[0] sky130_fd_sc_hd__conb_1
X_15181_ _08275_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__clkbuf_4
X_12393_ rbzero.tex_b1\[57\] rbzero.tex_b1\[56\] _04931_ vssd1 vssd1 vccd1 vccd1 _05578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__clkbuf_2
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ _04470_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19645__27 clknet_1_1__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
X_14063_ _07223_ _07232_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__nand2_1
X_18940_ _02481_ _02473_ _03052_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13014_ rbzero.wall_tracer.trackDistY\[-10\] _06188_ rbzero.wall_tracer.trackDistY\[-11\]
+ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__o211a_1
X_18871_ _03016_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17822_ _02108_ _02109_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__and2_1
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17753_ _01941_ _01948_ _01946_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a21o_1
X_14965_ _04437_ _04433_ _04438_ _04436_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__and4b_2
X_20558__18 clknet_1_0__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
XFILLER_82_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13916_ _06872_ _06867_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__and2b_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16704_ rbzero.traced_texa\[-2\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__a22o_1
X_17684_ _01862_ _01863_ _01754_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__or3b_1
XFILLER_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14896_ _08042_ _08035_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__nand2_1
X_19423_ _03335_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
X_16635_ _09601_ _09724_ vssd1 vssd1 vccd1 vccd1 _09725_ sky130_fd_sc_hd__xnor2_1
X_13847_ _06986_ _06988_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _09654_ _09655_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__nor2_1
X_19354_ rbzero.color_floor\[4\] _03290_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or2_1
X_13778_ _06742_ _06903_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__nand3b_1
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15517_ _08604_ _08611_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18305_ _02538_ _02539_ _02541_ _02542_ _04442_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o311a_1
X_12729_ _05891_ _05906_ net32 net33 vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and4b_1
X_19285_ rbzero.spi_registers.texadd3\[10\] _03255_ vssd1 vssd1 vccd1 vccd1 _03256_
+ sky130_fd_sc_hd__or2_1
X_16497_ _09480_ _09481_ _09586_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__nand3_1
XFILLER_176_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _02492_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__clkbuf_1
X_15448_ _08540_ _08542_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18167_ _02434_ _02435_ _02436_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__nor3_1
X_15379_ _08445_ _08471_ _08473_ _08455_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _10135_ _10136_ _10137_ _10131_ vssd1 vssd1 vccd1 vccd1 _10138_ sky130_fd_sc_hd__a211o_1
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18098_ _02376_ _02377_ _09852_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__o21ai_1
X_17049_ _09397_ _08497_ _09944_ _10069_ vssd1 vssd1 vccd1 vccd1 _10070_ sky130_fd_sc_hd__o31a_1
Xclkbuf_0__03787_ _03787_ vssd1 vssd1 vccd1 vccd1 clknet_0__03787_ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20060_ rbzero.debug_overlay.facingY\[-3\] _03658_ vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__or2_1
XFILLER_139_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ clknet_leaf_57_i_clk _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20306__171 clknet_1_1__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__inv_2
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20893_ clknet_leaf_53_i_clk _00482_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21514_ clknet_leaf_81_i_clk _01103_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21445_ net163 _01034_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21376_ clknet_leaf_7_i_clk _00965_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_162_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _04329_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20189_ _03761_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14750_ _06598_ _07917_ _06602_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__a21oi_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11962_ rbzero.debug_overlay.facingX\[-3\] _05110_ _05108_ rbzero.debug_overlay.facingX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a22o_1
XFILLER_85_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03776_ clknet_0__03776_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03776_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _06868_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__xnor2_1
X_10913_ _04252_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _07845_ _07851_ _07067_ _07332_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__and4b_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _05075_ _05081_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or2b_2
XFILLER_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16420_ _09485_ _09486_ _09510_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__a21o_1
X_13632_ _06797_ _06802_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__xor2_1
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10844_ _04216_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _09438_ _09439_ _09441_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__a21o_1
XFILLER_198_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13563_ _06730_ _06731_ _06732_ _06733_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__or4_1
X_10775_ rbzero.tex_g1\[15\] rbzero.tex_g1\[16\] _04177_ vssd1 vssd1 vccd1 vccd1 _04180_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15302_ _04464_ _08183_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__a21o_1
XFILLER_200_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19070_ rbzero.spi_registers.new_mapd\[5\] _03120_ _03131_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00774_ sky130_fd_sc_hd__o211a_1
X_12514_ _05382_ _05470_ _05551_ _05632_ _05646_ net7 vssd1 vssd1 vccd1 vccd1 _05696_
+ sky130_fd_sc_hd__mux4_1
X_16282_ _09008_ _09131_ _09372_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__o21ai_1
XFILLER_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13494_ _06618_ _06589_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nand2_1
X_18021_ _02237_ _02302_ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ _08313_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__buf_2
XFILLER_145_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ _04900_ _05553_ _05629_ _04702_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__o211a_1
XFILLER_200_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerY\[-5\] _08221_
+ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__or3_1
XFILLER_197_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12376_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _04978_ vssd1 vssd1 vccd1 vccd1 _05561_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14115_ _07213_ _07246_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__and2_1
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327_ rbzero.spi_registers.texadd1\[14\] vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__inv_2
X_19972_ _08241_ _03570_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nor2_1
X_15095_ rbzero.debug_overlay.playerY\[-8\] vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__inv_2
XFILLER_141_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14046_ _07196_ _07195_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__and2b_1
X_18923_ _03043_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11258_ _04449_ _03971_ _04446_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a21oi_1
XFILLER_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18854_ _03007_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11189_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _04395_ vssd1 vssd1 vccd1 vccd1 _04397_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17805_ _01842_ _02093_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__xor2_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15997_ _09089_ _09091_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__xor2_2
X_18785_ _02971_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17736_ _01937_ _01996_ _02024_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nand3_1
XFILLER_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ rbzero.wall_tracer.visualWallDist\[5\] _08046_ vssd1 vssd1 vccd1 vccd1 _08080_
+ sky130_fd_sc_hd__or2_1
XFILLER_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17667_ _01918_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__xnor2_1
X_14879_ rbzero.wall_tracer.stepDistY\[9\] _08029_ _07868_ vssd1 vssd1 vccd1 vccd1
+ _08030_ sky130_fd_sc_hd__mux2_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19406_ _03325_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
X_16618_ _09705_ _09707_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__nor2_1
XFILLER_165_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17598_ _01887_ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__nand2_1
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16549_ _09612_ _09613_ _09638_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__a21o_1
X_19337_ rbzero.color_sky\[3\] _03282_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or2_1
XFILLER_206_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19268_ rbzero.spi_registers.texadd3\[3\] _03242_ vssd1 vssd1 vccd1 vccd1 _03246_
+ sky130_fd_sc_hd__or2_1
XFILLER_206_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ rbzero.spi_registers.new_texadd\[2\]\[1\] _02481_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02482_ sky130_fd_sc_hd__mux2_1
X_19199_ rbzero.spi_registers.new_texadd\[1\]\[23\] _03173_ _03204_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__o211a_1
XFILLER_191_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21230_ clknet_leaf_11_i_clk _00819_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20336__197 clknet_1_1__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03808_ clknet_0__03808_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03808_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21161_ clknet_leaf_13_i_clk _00750_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20112_ rbzero.debug_overlay.vplaneY\[-2\] _03655_ _03710_ _03695_ vssd1 vssd1 vccd1
+ vccd1 _01237_ sky130_fd_sc_hd__a211o_1
XFILLER_131_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21092_ clknet_leaf_93_i_clk _00681_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20043_ rbzero.pov.ready_buffer\[42\] _03656_ _03672_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01206_ sky130_fd_sc_hd__o211a_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21994_ net140 _01583_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ clknet_leaf_51_i_clk _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_93_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20876_ clknet_leaf_68_i_clk _00465_ vssd1 vssd1 vccd1 vccd1 rbzero.side_hot sky130_fd_sc_hd__dfxtp_2
XFILLER_201_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ rbzero.tex_r0\[54\] rbzero.tex_r0\[53\] _04066_ vssd1 vssd1 vccd1 vccd1 _04067_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _04028_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12230_ rbzero.tex_g1\[24\] _04935_ _04933_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21428_ clknet_leaf_96_i_clk _01017_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _04932_ vssd1 vssd1 vccd1 vccd1 _05349_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_31_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_21359_ clknet_leaf_21_i_clk _00948_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _04356_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ _04652_ _04412_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nor2_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _08556_ _08557_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__nand2_1
X_11043_ _04320_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15851_ _08944_ _08945_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__xor2_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _07965_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__clkbuf_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15782_ _08875_ _08876_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__nor2_1
X_18570_ _02767_ _02770_ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ rbzero.wall_tracer.trackDistX\[4\] vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__inv_2
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17521_ _01811_ _01812_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__xor2_2
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _07900_ _07901_ _06577_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__mux2_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ rbzero.debug_overlay.vplaneY\[-2\] _05107_ _05113_ _05132_ _05133_ vssd1
+ vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a221o_1
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20441__292 clknet_1_1__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__inv_2
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _01742_ _01743_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__nand2_1
XFILLER_73_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14664_ _07409_ _07833_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__or2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ gpout0.hpos\[7\] _04639_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__nor2_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16403_ _09492_ _09493_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__nor2_1
X_13615_ _06722_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__nor2_1
X_10827_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _04203_ vssd1 vssd1 vccd1 vccd1 _04207_
+ sky130_fd_sc_hd__mux2_1
X_17383_ _08404_ _09076_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__or2_1
XFILLER_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14595_ _07755_ _07757_ _07762_ _07764_ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__o2111a_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19122_ rbzero.spi_registers.new_texadd\[0\]\[13\] _03155_ _03161_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__o211a_1
X_16334_ rbzero.wall_tracer.stepDistY\[8\] _08405_ _09190_ _09425_ vssd1 vssd1 vccd1
+ vccd1 _09426_ sky130_fd_sc_hd__a22o_2
XFILLER_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ _06657_ _06600_ _06713_ _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__o211ai_4
X_10758_ rbzero.tex_g1\[23\] rbzero.tex_g1\[24\] _04166_ vssd1 vssd1 vccd1 vccd1 _04171_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19053_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__clkbuf_2
XFILLER_199_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16265_ _09265_ _09266_ _09356_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__o21ai_1
X_13477_ _06512_ _06498_ _06603_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__mux2_1
X_10689_ _04134_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__clkbuf_1
X_18004_ _02216_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__xnor2_1
X_15216_ rbzero.wall_tracer.visualWallDist\[-2\] _08160_ vssd1 vssd1 vccd1 vccd1 _08311_
+ sky130_fd_sc_hd__or2_1
X_12428_ rbzero.tex_b1\[27\] _04926_ _04928_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__and3_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16196_ _09027_ _09170_ _09171_ _09172_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__a22o_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15147_ _08241_ rbzero.debug_overlay.playerY\[-5\] _06076_ vssd1 vssd1 vccd1 vccd1
+ _08242_ sky130_fd_sc_hd__mux2_1
X_12359_ _05047_ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__or2_1
XFILLER_181_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19955_ _03607_ _03609_ _03103_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__o21a_1
X_15078_ _07969_ _07970_ _08147_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ _07163_ _07164_ _07198_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__o21ai_1
X_18906_ rbzero.pov.spi_buffer\[60\] rbzero.pov.ready_buffer\[60\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19886_ _03555_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18837_ _02998_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20524__367 clknet_1_1__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__inv_2
X_18768_ _02929_ _02957_ rbzero.spi_registers.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1
+ _02960_ sky130_fd_sc_hd__a21oi_1
XFILLER_208_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17719_ _09662_ _02007_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__nor2_1
X_18699_ _02881_ _02884_ _02882_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a21bo_1
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20730_ _03935_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__buf_1
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20661_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03883_
+ sky130_fd_sc_hd__nand2_1
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20592_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03825_
+ sky130_fd_sc_hd__or2_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20418__272 clknet_1_1__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__inv_2
XFILLER_176_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21213_ clknet_leaf_7_i_clk _00802_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21144_ clknet_leaf_1_i_clk _00733_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21075_ clknet_leaf_81_i_clk _00664_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20026_ rbzero.debug_overlay.facingX\[-6\] _03658_ vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__or2_1
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ net503 _01566_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11730_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__buf_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ clknet_leaf_55_i_clk _00517_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ rbzero.row_render.size\[3\] _04837_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nand2_1
X_20859_ clknet_leaf_61_i_clk _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _06545_ _06558_ _06564_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__or3_1
X_10612_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _04088_ vssd1 vssd1 vccd1 vccd1 _04094_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ _07539_ _07548_ _07550_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__o21a_1
X_11592_ rbzero.traced_texVinit\[1\] rbzero.texV\[1\] rbzero.texV\[0\] rbzero.traced_texVinit\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__o211a_1
XFILLER_168_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ _06499_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__nand2_1
X_10543_ rbzero.tex_r0\[62\] rbzero.tex_r0\[61\] _04055_ vssd1 vssd1 vccd1 vccd1 _04058_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16050_ _09010_ _09019_ _09017_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__a21o_1
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19687__66 clknet_1_0__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13262_ rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__inv_2
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _04019_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15001_ _08110_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
X_12213_ _05393_ _05395_ _05397_ _05399_ _04967_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__o221a_1
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _04427_ _06046_ _06057_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__and3_1
XFILLER_123_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _04931_ vssd1 vssd1 vccd1 vccd1 _05332_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19740_ rbzero.pov.spi_buffer\[9\] rbzero.pov.spi_buffer\[10\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ _04832_ _05244_ _05262_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a31o_1
X_16952_ _09685_ _09566_ _09045_ vssd1 vssd1 vccd1 vccd1 _09974_ sky130_fd_sc_hd__a21o_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11026_ _04311_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
X_15903_ _08761_ _08764_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__nor2_1
XFILLER_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16883_ _09008_ _09363_ _09616_ _09904_ vssd1 vssd1 vccd1 vccd1 _09905_ sky130_fd_sc_hd__o31a_1
XFILLER_77_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18622_ _05132_ rbzero.debug_overlay.vplaneY\[-8\] vssd1 vssd1 vccd1 vccd1 _02827_
+ sky130_fd_sc_hd__nor2_1
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _08920_ _08926_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__xor2_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__or2_1
X_15765_ _08835_ _08858_ _08859_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__a21oi_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ rbzero.map_overlay.i_mapdy\[1\] _06089_ _06121_ rbzero.map_overlay.i_mapdy\[4\]
+ _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__a221o_1
XFILLER_205_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17504_ _01673_ _01682_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a21oi_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ _05082_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__nor2_4
X_14716_ _07884_ _07885_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__or2_1
X_15696_ _08734_ _08233_ _08484_ _08471_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__and4bb_1
X_18484_ _09866_ _06091_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__or3_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _09167_ _10093_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nor2_1
X_14647_ _06579_ _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__or2_1
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11859_ _04650_ _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__nor2_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 rbzero.spi_registers.vshift\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _10305_ _10381_ _10382_ vssd1 vssd1 vccd1 vccd1 _10384_ sky130_fd_sc_hd__and3_1
X_14578_ _07417_ _07444_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nor2_1
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ rbzero.spi_registers.new_texadd\[0\]\[6\] _03141_ _03151_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00789_ sky130_fd_sc_hd__o211a_1
X_16317_ _09290_ _09303_ _09304_ _09302_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__a22o_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13529_ _06633_ _06696_ _06699_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__a21o_2
X_17297_ _10315_ _08620_ _10313_ vssd1 vssd1 vccd1 vccd1 _10316_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16248_ _09338_ _09339_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__nand2_1
X_19036_ _08116_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__buf_6
XFILLER_103_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16179_ _08151_ _08731_ _08847_ _08166_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__o22ai_1
XFILLER_86_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19938_ _03594_ _03595_ _03561_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20448__298 clknet_1_1__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__inv_2
X_19869_ rbzero.pov.spi_buffer\[71\] rbzero.pov.spi_buffer\[72\] _03467_ vssd1 vssd1
+ vccd1 vccd1 _03547_ sky130_fd_sc_hd__mux2_1
XFILLER_29_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21900_ net426 _01489_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21831_ net357 _01420_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21762_ net288 _01351_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20713_ _03926_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21693_ net219 _01282_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20644_ _03865_ _03866_ _03860_ _03864_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__a211o_1
XFILLER_108_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20575_ _03811_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21127_ clknet_leaf_93_i_clk _00716_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21058_ clknet_leaf_97_i_clk _00647_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _06075_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__buf_4
X_20009_ rbzero.pov.ready_buffer\[57\] _03586_ _03649_ vssd1 vssd1 vccd1 vccd1 _03650_
+ sky130_fd_sc_hd__o21a_1
X_13880_ _06757_ _06729_ _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__a21oi_1
XFILLER_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and2_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15550_ _08641_ _08643_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__a21oi_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _05939_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _07580_ _07624_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__xor2_1
X_11713_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__buf_4
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _08503_ _08500_ _08501_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__a21o_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ net48 _05833_ _05846_ _05854_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a31o_1
XFILLER_15_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _10023_ _10115_ _10113_ vssd1 vssd1 vccd1 vccd1 _10240_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _07590_ _07594_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__xor2_1
XFILLER_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ _04819_ _04823_ _04825_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__or4_1
XFILLER_196_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03458_ clknet_0__03458_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03458_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17151_ _10160_ _10170_ vssd1 vssd1 vccd1 vccd1 _10171_ sky130_fd_sc_hd__xnor2_1
X_14363_ _07253_ _07248_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor2_1
XFILLER_195_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11575_ _04763_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__nor2_1
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_4
Xinput27 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_4
X_16102_ _08581_ _09053_ _09195_ _08461_ vssd1 vssd1 vccd1 vccd1 _09196_ sky130_fd_sc_hd__o22a_1
Xinput38 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_4
XFILLER_155_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13314_ _06474_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__and2_1
Xinput49 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_6
X_10526_ rbzero.tex_r1\[3\] rbzero.tex_r1\[4\] _04046_ vssd1 vssd1 vccd1 vccd1 _04047_
+ sky130_fd_sc_hd__mux2_1
X_17082_ _09968_ _09980_ vssd1 vssd1 vccd1 vccd1 _10103_ sky130_fd_sc_hd__or2_1
XFILLER_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _07462_ _07464_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__or2b_1
XFILLER_156_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _09023_ _09001_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__or2b_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13245_ _06324_ _06328_ _06331_ _06322_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__a31o_1
XFILLER_196_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10457_ _04010_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13176_ _06305_ _06307_ _06308_ _06295_ _06292_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a32o_1
X_10388_ gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__buf_4
XFILLER_112_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _05314_ vssd1 vssd1 vccd1 vccd1 _05315_
+ sky130_fd_sc_hd__mux2_1
XFILLER_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17984_ _02088_ _02253_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__or2b_1
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19723_ rbzero.pov.spi_buffer\[1\] rbzero.pov.spi_buffer\[2\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16935_ _09670_ _09184_ _08516_ vssd1 vssd1 vccd1 vccd1 _09957_ sky130_fd_sc_hd__a21oi_1
X_12058_ rbzero.tex_r1\[61\] _05199_ _05032_ _04890_ vssd1 vssd1 vccd1 vccd1 _05247_
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11009_ _04302_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
X_16866_ rbzero.wall_tracer.trackDistX\[-1\] _09888_ _09844_ vssd1 vssd1 vccd1 vccd1
+ _09889_ sky130_fd_sc_hd__mux2_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18605_ _02794_ rbzero.wall_tracer.rayAddendY\[0\] _02797_ vssd1 vssd1 vccd1 vccd1
+ _02811_ sky130_fd_sc_hd__o21a_1
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15817_ _08213_ _08343_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__nor2_1
X_19585_ _03421_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16797_ _09817_ _09818_ _09819_ vssd1 vssd1 vccd1 vccd1 _09827_ sky130_fd_sc_hd__a21bo_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18536_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__nor2_1
X_15748_ _08252_ _08440_ _08791_ _08790_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__or4b_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _02690_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15679_ _08246_ _08337_ _08343_ _08265_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__o22a_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17418_ _01704_ _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__nand2_1
X_20300__166 clknet_1_1__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__inv_2
X_18398_ _02616_ _02621_ _02628_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__o21ai_1
XFILLER_14_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17349_ _10366_ _10367_ vssd1 vssd1 vccd1 vccd1 _10368_ sky130_fd_sc_hd__nand2_1
XFILLER_14_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ _05644_ _09728_ _03092_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__and3_1
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22030_ clknet_leaf_54_i_clk _01619_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20229__101 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__inv_2
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20381__238 clknet_1_1__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__inv_2
XFILLER_29_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21814_ net340 _01403_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21745_ net271 _01334_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21676_ clknet_leaf_0_i_clk _01265_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20275__143 clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__inv_2
XFILLER_196_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20627_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03854_
+ sky130_fd_sc_hd__or2_1
XFILLER_32_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ rbzero.spi_registers.texadd0\[21\] _04535_ _04551_ vssd1 vssd1 vccd1 vccd1
+ _04552_ sky130_fd_sc_hd__o21ai_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ rbzero.spi_registers.texadd3\[9\] _04465_ _04456_ rbzero.spi_registers.texadd2\[9\]
+ _04470_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a221o_1
XFILLER_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13030_ rbzero.wall_tracer.trackDistY\[2\] _06172_ _06202_ rbzero.wall_tracer.trackDistY\[1\]
+ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__o221a_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14981_ rbzero.wall_tracer.stepDistX\[-4\] _07964_ _08092_ vssd1 vssd1 vccd1 vccd1
+ _08100_ sky130_fd_sc_hd__mux2_1
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16720_ _04437_ _04433_ _05050_ _09729_ vssd1 vssd1 vccd1 vccd1 _09760_ sky130_fd_sc_hd__nand4_4
X_13932_ _06782_ _06887_ _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__o21a_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13863_ _06951_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__xnor2_1
X_16651_ _04638_ _05079_ _09732_ vssd1 vssd1 vccd1 vccd1 _09736_ sky130_fd_sc_hd__and3_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15602_ _08327_ _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__nor2_1
X_12814_ _05988_ _05942_ _05990_ _05946_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a22o_2
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19370_ rbzero.spi_registers.new_vshift\[4\] _03297_ _03304_ _03302_ vssd1 vssd1
+ vccd1 vccd1 _00901_ sky130_fd_sc_hd__o211a_1
X_16582_ _08434_ _09669_ _09671_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__o21ba_1
X_13794_ _06914_ _06915_ _06921_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__or3_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18321_ _09749_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__buf_6
X_15533_ _08614_ _08627_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__xnor2_1
X_12745_ net46 _05920_ _05921_ net43 _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a221o_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15464_ _08556_ _08557_ _08558_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__a21o_1
XFILLER_176_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18252_ rbzero.spi_registers.new_texadd\[2\]\[15\] rbzero.spi_registers.spi_buffer\[15\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ net46 _05843_ _05846_ _05854_ net43 vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a32o_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17203_ _10220_ _10222_ vssd1 vssd1 vccd1 vccd1 _10223_ sky130_fd_sc_hd__xor2_1
XFILLER_175_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14415_ _07584_ _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__nand2_1
XFILLER_169_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__buf_4
X_15395_ _08487_ _08489_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__and2_1
X_18183_ _02449_ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nor2_1
XFILLER_184_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17134_ _10151_ _10152_ vssd1 vssd1 vccd1 vccd1 _10154_ sky130_fd_sc_hd__or2_1
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14346_ _07515_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__nor2_1
XFILLER_200_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ _04746_ _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__and2_1
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17065_ _10081_ _10085_ vssd1 vssd1 vccd1 vccd1 _10086_ sky130_fd_sc_hd__xnor2_1
X_10509_ rbzero.tex_r1\[11\] rbzero.tex_r1\[12\] _04035_ vssd1 vssd1 vccd1 vccd1 _04038_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14277_ _06720_ _07209_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__nor2_1
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11489_ rbzero.debug_overlay.playerX\[0\] vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__inv_2
XFILLER_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _08994_ _08996_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__xor2_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ rbzero.wall_tracer.visualWallDist\[0\] _06327_ _04443_ vssd1 vssd1 vccd1
+ vccd1 _06399_ sky130_fd_sc_hd__a21o_1
XFILLER_48_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _06322_ _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XFILLER_98_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _02184_ _02185_ _02254_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a21o_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16918_ _09938_ _09939_ vssd1 vssd1 vccd1 vccd1 _09940_ sky130_fd_sc_hd__and2_1
XFILLER_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17898_ _02091_ _02094_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__and2_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19637_ _03453_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16849_ _09872_ _09593_ vssd1 vssd1 vccd1 vccd1 _09873_ sky130_fd_sc_hd__nand2_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19568_ _03412_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18519_ rbzero.debug_overlay.playerX\[3\] _02733_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _02734_ sky130_fd_sc_hd__mux2_1
XFILLER_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ _03376_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21530_ clknet_leaf_97_i_clk _01119_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21461_ net179 _01050_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20412_ clknet_1_0__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__buf_1
XFILLER_175_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21392_ clknet_leaf_11_i_clk _00981_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22013_ clknet_leaf_68_i_clk _01602_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03792_ clknet_0__03792_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03792_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10860_ _04224_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _04143_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__buf_4
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ net54 vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__clkbuf_8
XFILLER_185_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21728_ net254 _01317_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ net5 vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__inv_2
XFILLER_185_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21659_ clknet_leaf_17_i_clk _01248_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _07367_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
X_11412_ _04496_ _04497_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__nand2_1
X_15180_ _08269_ _08274_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__or2_1
X_12392_ _05575_ _05576_ _05190_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_83 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_83/HI o_rgb[10] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_94 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_94/HI zeros[1] sky130_fd_sc_hd__conb_1
XFILLER_166_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ _07254_ _07285_ _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__o21ai_2
XFILLER_158_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ _04467_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_67_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14062_ _07223_ _07232_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or2_1
X_11274_ _04465_ rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__nand2_1
XFILLER_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13013_ rbzero.wall_tracer.trackDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__inv_2
X_18870_ rbzero.pov.spi_buffer\[43\] rbzero.pov.ready_buffer\[43\] _03011_ vssd1 vssd1
+ vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17821_ _02108_ _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__nor2_1
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ _01927_ _01935_ _01933_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a21o_1
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14964_ rbzero.wall_tracer.visualWallDist\[10\] _08047_ _08090_ _08085_ vssd1 vssd1
+ vccd1 vccd1 _00434_ sky130_fd_sc_hd__o211a_1
XFILLER_75_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16703_ rbzero.traced_texa\[-3\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22o_1
X_13915_ _07065_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17683_ _01972_ _01973_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__nand2_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14895_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _08042_
+ sky130_fd_sc_hd__inv_2
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19422_ _02489_ rbzero.spi_registers.new_leak\[5\] _03329_ vssd1 vssd1 vccd1 vccd1
+ _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16634_ _09721_ _09723_ vssd1 vssd1 vccd1 vccd1 _09724_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ _07001_ _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__nand2_1
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19353_ rbzero.color_floor\[3\] _03289_ _03294_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__a21o_1
X_16565_ _09393_ _09529_ _09531_ _09532_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__a22oi_2
X_13777_ _06729_ _06758_ _06901_ _06902_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__a22o_1
X_10989_ _04143_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18304_ _02538_ _02539_ _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o21ai_1
X_15516_ _08609_ _08610_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__nand2_1
XFILLER_149_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ _05899_ _05900_ _05903_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a22o_1
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19284_ _03241_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__buf_2
XFILLER_206_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16496_ _09480_ _09481_ _09586_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__a21o_2
XFILLER_15_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18235_ rbzero.spi_registers.new_texadd\[2\]\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _02479_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
X_15447_ _08171_ _08541_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__or2_1
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12659_ _05829_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__or2_1
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] _02431_
+ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ _08472_ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__buf_2
XFILLER_156_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _10128_ vssd1 vssd1 vccd1 vccd1 _10137_ sky130_fd_sc_hd__inv_2
X_14329_ _07488_ _07494_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__xor2_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18097_ _02374_ _02375_ _09866_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a21o_1
XFILLER_143_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03786_ _03786_ vssd1 vssd1 vccd1 vccd1 clknet_0__03786_ sky130_fd_sc_hd__clkbuf_16
X_17048_ _09941_ _09942_ vssd1 vssd1 vccd1 vccd1 _10069_ sky130_fd_sc_hd__nand2_1
XFILLER_143_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18999_ rbzero.spi_registers.mosi rbzero.spi_registers.mosi_buffer\[0\] _03084_ vssd1
+ vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20961_ clknet_leaf_57_i_clk _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20892_ clknet_leaf_44_i_clk _00481_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20493__339 clknet_1_0__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__inv_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21513_ clknet_leaf_81_i_clk _01102_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21444_ net162 _01033_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21375_ clknet_leaf_24_i_clk _00964_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20387__244 clknet_1_0__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__inv_2
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20257_ clknet_1_1__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__buf_1
XFILLER_27_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20188_ rbzero.spi_registers.new_texadd\[3\]\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__mux2_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ rbzero.debug_overlay.facingX\[-2\] _05107_ _05113_ rbzero.debug_overlay.facingX\[-4\]
+ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a221o_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10912_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _04248_ vssd1 vssd1 vccd1 vccd1 _04252_
+ sky130_fd_sc_hd__mux2_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _06869_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__xnor2_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _07206_ _07398_ _07337_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__o21ba_1
XFILLER_189_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11892_ _04638_ _05079_ _05078_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__a21oi_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ _06748_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__xnor2_1
X_10843_ rbzero.tex_g0\[48\] rbzero.tex_g0\[47\] _04215_ vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _09438_ _09439_ _09441_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__nand3_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13562_ _06701_ _06702_ _06703_ _06706_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__o211a_2
XFILLER_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10774_ _04179_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15301_ _08395_ _06044_ _06045_ _08147_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__a31o_1
X_12513_ _05646_ _05297_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__nand2_1
X_16281_ _08335_ _09131_ _09372_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__or3_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13493_ _06521_ _06590_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__nor2_1
XFILLER_160_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ _02303_ _02306_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__xnor2_1
X_15232_ _08325_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__clkbuf_4
X_12444_ _04900_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__nand2_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ rbzero.debug_overlay.playerY\[-4\] vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__inv_2
X_12375_ _05558_ _05559_ _05190_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__mux2_1
XFILLER_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _07256_ _07284_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__xnor2_4
XFILLER_197_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ rbzero.spi_registers.texadd0\[14\] _04467_ vssd1 vssd1 vccd1 vccd1 _04518_
+ sky130_fd_sc_hd__or2_1
XFILLER_180_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19971_ _03611_ _03620_ _03621_ _03579_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__o211a_1
X_15094_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18922_ rbzero.pov.spi_buffer\[68\] rbzero.pov.ready_buffer\[68\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
X_14045_ _07168_ _07192_ _07193_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__and3_1
XFILLER_140_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11257_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__inv_4
XFILLER_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18853_ rbzero.pov.spi_buffer\[35\] rbzero.pov.ready_buffer\[35\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
X_11188_ _04396_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17804_ _02033_ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__xor2_2
XFILLER_209_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18784_ rbzero.pov.spi_buffer\[2\] rbzero.pov.ready_buffer\[2\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15996_ _08614_ _08627_ _09090_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__a21oi_2
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17735_ _01937_ _01996_ _02024_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a21o_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.trackDistX\[5\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__mux2_1
XFILLER_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17666_ _01955_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__xor2_1
X_14878_ _06600_ _07995_ _07866_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__o21ai_2
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19405_ _02489_ rbzero.spi_registers.new_floor\[5\] _03319_ vssd1 vssd1 vccd1 vccd1
+ _03325_ sky130_fd_sc_hd__mux2_1
X_16617_ _09541_ _09577_ _09706_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ _06991_ _06980_ _06989_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__nor3_1
X_17597_ _01885_ _01886_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__or2_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19336_ rbzero.color_sky\[2\] _03280_ _03284_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__a21o_1
X_16548_ _09623_ _09637_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19267_ rbzero.spi_registers.new_texadd\[3\]\[2\] _03240_ _03245_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00857_ sky130_fd_sc_hd__o211a_1
X_16479_ _09427_ _09430_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__nand2_1
XFILLER_164_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18218_ rbzero.spi_registers.spi_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__buf_4
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19198_ rbzero.spi_registers.texadd1\[23\] _03175_ vssd1 vssd1 vccd1 vccd1 _03204_
+ sky130_fd_sc_hd__or2_1
XFILLER_15_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03807_ clknet_0__03807_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03807_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18149_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21160_ clknet_leaf_13_i_clk _00749_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20111_ rbzero.pov.ready_buffer\[7\] _03687_ _03664_ vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__and3_1
XFILLER_160_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21091_ clknet_leaf_97_i_clk _00680_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20042_ rbzero.debug_overlay.facingX\[0\] _03658_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__or2_1
XFILLER_59_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21993_ net139 _01582_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20944_ clknet_leaf_52_i_clk _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ clknet_leaf_20_i_clk _00464_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_hot\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_183_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ rbzero.tex_r1\[20\] rbzero.tex_r1\[21\] _04024_ vssd1 vssd1 vccd1 vccd1 _04028_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21427_ clknet_leaf_96_i_clk _01016_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_19702__79 clknet_1_0__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
XFILLER_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12160_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _05002_ vssd1 vssd1 vccd1 vccd1 _05348_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21358_ clknet_leaf_21_i_clk _00947_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11111_ rbzero.tex_b0\[48\] rbzero.tex_b0\[47\] _04351_ vssd1 vssd1 vccd1 vccd1 _04356_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ _04654_ _04655_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nand2_1
X_21289_ clknet_leaf_6_i_clk _00878_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ rbzero.tex_b1\[16\] rbzero.tex_b1\[17\] _04314_ vssd1 vssd1 vccd1 vccd1 _04320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _08304_ _08458_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__nor2_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801_ rbzero.wall_tracer.stepDistY\[-4\] _07964_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07965_ sky130_fd_sc_hd__mux2_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _08847_ _08473_ _08458_ _08274_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__o22a_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ rbzero.wall_tracer.trackDistX\[5\] vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__inv_2
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ rbzero.wall_tracer.visualWallDist\[3\] _08475_ _08445_ vssd1 vssd1 vccd1
+ vccd1 _01812_ sky130_fd_sc_hd__and3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _07806_ _07805_ _07810_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__a21o_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ rbzero.debug_overlay.vplaneY\[-5\] _05112_ _04652_ vssd1 vssd1 vccd1 vccd1
+ _05133_ sky130_fd_sc_hd__a21bo_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17451_ _01742_ _01743_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nor2_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ _04656_ _04655_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nor2_2
X_14663_ _07409_ _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__nand2_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _08616_ _09491_ _09489_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__o21a_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10826_ _04206_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__clkbuf_1
X_13614_ _06682_ _06784_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__nand2_2
X_17382_ _01674_ _10314_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__nand2_1
XFILLER_60_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14594_ _06982_ _07159_ _07758_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__and3b_1
XFILLER_164_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19121_ rbzero.spi_registers.texadd0\[13\] _03156_ vssd1 vssd1 vccd1 vccd1 _03161_
+ sky130_fd_sc_hd__or2_1
XFILLER_201_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16333_ _09423_ _09308_ _09424_ _08144_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__a211o_1
XFILLER_199_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10757_ _04170_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13545_ _06595_ _06714_ _06715_ _06581_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__a211o_1
XFILLER_185_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19052_ rbzero.spi_registers.got_new_mapd _03100_ vssd1 vssd1 vccd1 vccd1 _03121_
+ sky130_fd_sc_hd__and2_1
X_16264_ _09162_ _09240_ _09264_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__a21o_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _06569_ _06538_ _06554_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and3_1
X_10688_ rbzero.tex_g1\[56\] rbzero.tex_g1\[57\] _04132_ vssd1 vssd1 vccd1 vccd1 _04134_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003_ _08455_ _09243_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__nor2_1
XFILLER_139_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12427_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _04893_ vssd1 vssd1 vccd1 vccd1 _05612_
+ sky130_fd_sc_hd__mux2_1
X_15215_ _08309_ rbzero.debug_overlay.playerY\[-2\] _06076_ vssd1 vssd1 vccd1 vccd1
+ _08310_ sky130_fd_sc_hd__mux2_1
X_16195_ _09268_ _09287_ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _05472_ _05543_ _04899_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__mux2_1
X_15146_ rbzero.debug_overlay.playerY\[-5\] _08221_ vssd1 vssd1 vccd1 vccd1 _08241_
+ sky130_fd_sc_hd__xor2_1
XFILLER_141_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11309_ rbzero.texu_hot\[2\] _04488_ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15077_ _08152_ _08164_ _08166_ _08171_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__or4_2
X_19954_ rbzero.pov.ready_buffer\[73\] _03586_ _03569_ _03608_ vssd1 vssd1 vccd1 vccd1
+ _03609_ sky130_fd_sc_hd__o211a_1
XFILLER_99_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12289_ _05473_ _05474_ _04946_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__mux2_1
XFILLER_45_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14028_ _07163_ _07164_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__or3_1
X_18905_ _03034_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19885_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] _08116_ vssd1 vssd1
+ vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18836_ rbzero.pov.spi_buffer\[27\] rbzero.pov.ready_buffer\[27\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18767_ rbzero.spi_registers.spi_counter\[4\] _02929_ _02957_ vssd1 vssd1 vccd1 vccd1
+ _02959_ sky130_fd_sc_hd__and3_1
X_15979_ _08570_ _08546_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__or2b_1
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ _09662_ _02007_ _01901_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__or3_1
X_18698_ rbzero.debug_overlay.vplaneY\[-1\] _02879_ vssd1 vssd1 vccd1 vccd1 _02898_
+ sky130_fd_sc_hd__nand2_1
XFILLER_63_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17649_ _01919_ _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20660_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03882_
+ sky130_fd_sc_hd__or2_1
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19319_ rbzero.spi_registers.new_leak\[1\] _03271_ _03274_ _03265_ vssd1 vssd1 vccd1
+ vccd1 _00880_ sky130_fd_sc_hd__o211a_1
XFILLER_91_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20591_ rbzero.texV\[-9\] _03695_ _03819_ _03824_ vssd1 vssd1 vccd1 vccd1 _01602_
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21212_ clknet_leaf_5_i_clk _00801_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21143_ clknet_leaf_1_i_clk _00732_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21074_ clknet_leaf_81_i_clk _00663_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20025_ rbzero.pov.ready_buffer\[35\] _03656_ _03661_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01199_ sky130_fd_sc_hd__o211a_1
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20499__345 clknet_1_0__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__inv_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ net502 _01565_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ clknet_leaf_55_i_clk _00516_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ rbzero.row_render.size\[4\] _04838_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20858_ clknet_leaf_62_i_clk _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _04093_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11591_ rbzero.texV\[3\] _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__xor2_2
XFILLER_70_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20789_ _03965_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__clkbuf_1
X_13330_ _06377_ _06500_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__xor2_4
X_10542_ _04057_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13261_ _06431_ _06424_ _06428_ _06411_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__a211o_1
X_10473_ rbzero.tex_r1\[28\] rbzero.tex_r1\[29\] _04013_ vssd1 vssd1 vccd1 vccd1 _04019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12212_ rbzero.tex_g1\[0\] _04935_ _04933_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_
+ sky130_fd_sc_hd__a31o_1
X_15000_ rbzero.wall_tracer.stepDistX\[5\] _08015_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08110_ sky130_fd_sc_hd__mux2_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13192_ rbzero.wall_tracer.visualWallDist\[-5\] _06327_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a21o_1
XFILLER_136_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _04932_ vssd1 vssd1 vccd1 vccd1 _05331_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12074_ net42 vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__buf_6
X_16951_ _09970_ _09972_ _08950_ vssd1 vssd1 vccd1 vccd1 _09973_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ rbzero.tex_b1\[24\] rbzero.tex_b1\[25\] _04303_ vssd1 vssd1 vccd1 vccd1 _04311_
+ sky130_fd_sc_hd__mux2_1
X_15902_ _08763_ _08811_ _08994_ _08996_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__a2bb2o_2
X_16882_ _09498_ _09615_ vssd1 vssd1 vccd1 vccd1 _09904_ sky130_fd_sc_hd__nand2_1
XFILLER_106_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18621_ rbzero.debug_overlay.vplaneY\[-2\] _05129_ vssd1 vssd1 vccd1 vccd1 _02826_
+ sky130_fd_sc_hd__xor2_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _08914_ _08927_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__and2_1
XFILLER_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _02761_ _02762_ _08136_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _08799_ _08836_ _08857_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__and3_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ rbzero.map_overlay.i_mapdy\[2\] rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1
+ _06152_ sky130_fd_sc_hd__xor2_1
XFILLER_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17503_ _01674_ _10314_ _01681_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a21oi_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _06613_ _07817_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__nor2_1
XFILLER_205_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11927_ _05073_ _05089_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__or2_4
X_18483_ _06088_ _06090_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__nor2_1
XFILLER_79_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15695_ _08734_ _08473_ _08457_ _08233_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__o22ai_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _10096_ _10344_ _10221_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a21o_1
XFILLER_127_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14646_ _07793_ _07795_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__xnor2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _04703_ _04745_ _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__o22a_1
XFILLER_199_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17365_ _10305_ _10381_ _10382_ vssd1 vssd1 vccd1 vccd1 _10383_ sky130_fd_sc_hd__a21oi_2
X_10809_ _04197_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_19 rbzero.spi_registers.vshift\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11789_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _04978_ vssd1 vssd1 vccd1 vccd1 _04979_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14577_ _07640_ _07722_ _07740_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__o21a_1
X_19104_ rbzero.spi_registers.texadd0\[6\] _03143_ vssd1 vssd1 vccd1 vccd1 _03151_
+ sky130_fd_sc_hd__or2_1
X_16316_ _09406_ _08409_ _09294_ _09407_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__o31ai_1
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13528_ _06595_ _06656_ _06698_ _06655_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__o211a_1
X_17296_ _08399_ vssd1 vssd1 vccd1 vccd1 _10315_ sky130_fd_sc_hd__buf_2
XFILLER_173_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19035_ rbzero.map_overlay.i_othery\[1\] _03101_ vssd1 vssd1 vccd1 vccd1 _03109_
+ sky130_fd_sc_hd__or2_1
X_16247_ _09338_ _09339_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__or2_2
XFILLER_185_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13459_ _06566_ _06572_ _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16178_ _08151_ _08165_ _08731_ _08847_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__or4_1
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _06034_ _06074_ _08223_ _08157_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__a31o_1
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19937_ _04674_ _03591_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__or2_1
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19868_ _03546_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18819_ _02967_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__clkbuf_4
X_19799_ _03510_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21830_ net356 _01419_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21761_ net287 _01350_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20712_ _04442_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__and2_1
XFILLER_169_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21692_ net218 _01281_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20643_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__inv_2
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20574_ _03728_ _03809_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_45_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19692__70 clknet_1_0__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21126_ clknet_leaf_92_i_clk _00715_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21057_ clknet_leaf_99_i_clk _00646_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20507__352 clknet_1_1__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__inv_2
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20008_ _03556_ _03648_ _03616_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__o21a_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12830_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nor2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ reg_gpout\[4\] clknet_1_1__leaf__05938_ net45 vssd1 vssd1 vccd1 vccd1 _05939_
+ sky130_fd_sc_hd__mux2_2
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ net485 _01548_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _07628_ _07670_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__nor2_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _04812_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__buf_6
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _08503_ _08500_ _08501_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__nand3_1
X_12692_ net52 _05842_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a21o_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11643_ _04827_ _04831_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__or3_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _07556_ _07567_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03457_ clknet_0__03457_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03457_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17150_ _10168_ _10169_ vssd1 vssd1 vccd1 vccd1 _10170_ sky130_fd_sc_hd__nor2_1
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11574_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _04764_ sky130_fd_sc_hd__nor2_1
X_14362_ _07532_ _07253_ _07309_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__or3b_1
XFILLER_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_6
XFILLER_195_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_4
X_16101_ _09194_ _09191_ _09045_ vssd1 vssd1 vccd1 vccd1 _09195_ sky130_fd_sc_hd__a21o_4
XFILLER_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_4
X_10525_ _03979_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13313_ _06448_ _06467_ _06477_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__and4_1
X_17081_ _09968_ _09980_ vssd1 vssd1 vccd1 vccd1 _10102_ sky130_fd_sc_hd__nand2_1
XFILLER_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14293_ _07455_ _07456_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__o21ai_2
XFILLER_196_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20252__122 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__inv_2
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16032_ _09093_ _09095_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__or2_2
X_13244_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__clkbuf_4
X_10456_ rbzero.tex_r1\[36\] rbzero.tex_r1\[37\] _04002_ vssd1 vssd1 vccd1 vccd1 _04010_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13175_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__nand2_1
XFILLER_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _04913_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__buf_4
XFILLER_124_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17983_ _02169_ _02255_ _02257_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a21o_1
XFILLER_105_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19722_ _03470_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
X_16934_ _09679_ _09681_ _09682_ _09678_ vssd1 vssd1 vccd1 vccd1 _09956_ sky130_fd_sc_hd__a2bb2o_1
X_12057_ rbzero.tex_r1\[63\] _05002_ _05245_ _04922_ vssd1 vssd1 vccd1 vccd1 _05246_
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11008_ rbzero.tex_b1\[32\] rbzero.tex_b1\[33\] _04292_ vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16865_ _09885_ _09886_ _09887_ vssd1 vssd1 vccd1 vccd1 _09888_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or2_1
X_15816_ _08195_ _08337_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__or2_1
XFILLER_93_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19584_ rbzero.spi_registers.new_texadd\[1\]\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__mux2_1
X_16796_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09826_ sky130_fd_sc_hd__nand2_1
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__nand2_1
XFILLER_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15747_ _08840_ _08793_ _08786_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__a21o_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12959_ rbzero.debug_overlay.playerX\[4\] _06129_ _06130_ rbzero.debug_overlay.playerY\[0\]
+ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__a221o_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18466_ _02667_ _02677_ _02691_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__o21ai_1
X_15678_ _08771_ _08772_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__or2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17417_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__xor2_1
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14629_ _07524_ _07579_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__nor2_1
X_18397_ _02569_ rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _02628_
+ sky130_fd_sc_hd__xor2_1
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17348_ _10144_ _10365_ vssd1 vssd1 vccd1 vccd1 _10367_ sky130_fd_sc_hd__or2_1
XFILLER_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17279_ _10296_ _10297_ vssd1 vssd1 vccd1 vccd1 _10298_ sky130_fd_sc_hd__nor2_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19018_ rbzero.spi_registers.got_new_other _03097_ vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__nand2_4
X_20290_ clknet_1_1__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__buf_1
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21813_ net339 _01402_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21744_ net270 _01333_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21675_ clknet_leaf_100_i_clk _01264_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20626_ rbzero.texV\[-3\] _03814_ _03819_ _03853_ vssd1 vssd1 vccd1 vccd1 _01608_
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11290_ rbzero.spi_registers.texadd1\[9\] _04460_ vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__and2_1
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21109_ clknet_leaf_92_i_clk _00698_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_14980_ _08099_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13931_ _06850_ _06886_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__nand2_1
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ net63 _05061_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__nor2_1
X_13862_ _06757_ _06728_ _07019_ _07032_ _07022_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__a32o_1
XFILLER_41_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15601_ _08358_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__buf_2
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ _05949_ net39 _05977_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__and4_1
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16581_ _09670_ _09184_ _08889_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13793_ _06914_ _06915_ _06921_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ rbzero.wall_tracer.rayAddendX\[-2\] _02527_ _02553_ _02556_ vssd1 vssd1 vccd1
+ vccd1 _00599_ sky130_fd_sc_hd__o22a_1
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15532_ _08625_ _08626_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__nor2_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12744_ net31 net30 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__or2_1
XFILLER_128_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18251_ _02500_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _08235_ _08328_ _08325_ _08253_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__o22a_1
XFILLER_163_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05842_ _05846_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__and2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17202_ _10091_ _10096_ _10221_ vssd1 vssd1 vccd1 vccd1 _10222_ sky130_fd_sc_hd__a21o_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14414_ _06942_ _07209_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__nor2_1
X_11626_ _04786_ _04806_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__or3b_1
X_18182_ _02440_ _02442_ _02441_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__o21ba_1
X_15394_ _08400_ _08440_ _08487_ _08488_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__or4bb_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _10151_ _10152_ vssd1 vssd1 vccd1 vccd1 _10153_ sky130_fd_sc_hd__nand2_1
XFILLER_184_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14345_ _07499_ _07514_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__and2_1
XFILLER_183_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11557_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _04747_
+ sky130_fd_sc_hd__or2_1
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _10083_ _10084_ vssd1 vssd1 vccd1 vccd1 _10085_ sky130_fd_sc_hd__xnor2_1
X_10508_ _04037_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14276_ _07210_ _07362_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__nand2_1
X_11488_ _04670_ rbzero.debug_overlay.playerY\[4\] rbzero.debug_overlay.playerX\[1\]
+ _04414_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__o221a_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16015_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerX\[-8\] _04464_
+ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__mux2_1
X_10439_ rbzero.tex_r1\[44\] rbzero.tex_r1\[45\] _03991_ vssd1 vssd1 vccd1 vccd1 _04001_
+ sky130_fd_sc_hd__mux2_1
X_13227_ _06396_ _06397_ _04444_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ rbzero.wall_tracer.visualWallDist\[5\] _04428_ _06324_ _06328_ vssd1 vssd1
+ vccd1 vccd1 _06329_ sky130_fd_sc_hd__o211a_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19671__51 clknet_1_0__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_12109_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__inv_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _02088_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__xor2_1
X_13089_ _06161_ _06258_ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__o21ai_4
XFILLER_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16917_ _09519_ _08620_ _09937_ vssd1 vssd1 vccd1 vccd1 _09939_ sky130_fd_sc_hd__o21ai_1
X_17897_ _01992_ _02166_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__nand2_1
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16848_ _06104_ vssd1 vssd1 vccd1 vccd1 _09872_ sky130_fd_sc_hd__buf_4
X_19636_ _03451_ _03440_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__and3b_1
XFILLER_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19567_ rbzero.spi_registers.new_texadd\[1\]\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
X_16779_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ _09808_ _09809_ vssd1 vssd1 vccd1 vccd1 _09811_ sky130_fd_sc_hd__a22oi_1
X_18518_ _09772_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19498_ rbzero.spi_registers.new_mapd\[13\] rbzero.spi_registers.spi_buffer\[13\]
+ _03361_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20259__128 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__inv_2
X_18449_ _09753_ _02666_ _02667_ _02676_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a31o_1
XFILLER_178_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21460_ net178 _01049_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21391_ clknet_leaf_10_i_clk _00980_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22012_ clknet_leaf_50_i_clk _01601_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03791_ clknet_0__03791_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03791_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10790_ _04187_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21727_ net253 _01316_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21658_ clknet_leaf_17_i_clk _01247_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_1
X_12460_ net8 _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__nand2_1
X_20470__318 clknet_1_0__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__inv_2
XFILLER_184_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _04496_ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__and2_1
X_12391_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _04931_ vssd1 vssd1 vccd1 vccd1 _05576_
+ sky130_fd_sc_hd__mux2_1
X_20609_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03839_
+ sky130_fd_sc_hd__nand2_1
Xtop_ew_algofoogle_84 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_84/HI o_rgb[11] sky130_fd_sc_hd__conb_1
X_21589_ clknet_leaf_16_i_clk _01178_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\]
+ sky130_fd_sc_hd__dfxtp_2
Xtop_ew_algofoogle_95 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_95/HI zeros[2] sky130_fd_sc_hd__conb_1
XFILLER_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _07286_ _07284_ _07298_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__a211o_1
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11342_ _04530_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__and2_1
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ _07187_ _07231_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__xnor2_1
X_11273_ _04459_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13012_ rbzero.wall_tracer.trackDistX\[-10\] vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__inv_2
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17820_ _01818_ _09560_ _02051_ _02050_ _01928_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__o32a_1
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20364__223 clknet_1_0__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__inv_2
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _02039_ _02040_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__nor2_1
X_14963_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.trackDistY\[10\] _08035_
+ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__a21o_1
XFILLER_102_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16702_ rbzero.traced_texa\[-4\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13914_ _07073_ _07084_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__xor2_2
XFILLER_43_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17682_ _01970_ _01971_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__nand2_1
XFILLER_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14894_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.trackDistX\[-10\]
+ _08037_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__mux2_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19421_ _03334_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
X_16633_ _09121_ _09722_ vssd1 vssd1 vccd1 vccd1 _09723_ sky130_fd_sc_hd__xnor2_1
X_13845_ _06992_ _07000_ _06999_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__o21ai_1
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19352_ rbzero.spi_registers.new_floor\[3\] rbzero.spi_registers.got_new_floor _03097_
+ _04409_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a31o_1
X_16564_ _09529_ _09653_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13776_ _06932_ _06945_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10988_ _04291_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18303_ _02540_ _02530_ _02529_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a21oi_1
X_15515_ _08605_ _08606_ _08608_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__nand3_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _05889_ _05904_ _05888_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__o21a_1
X_19283_ _03239_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__clkbuf_4
X_16495_ _09483_ _09585_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19708__85 clknet_1_1__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
XFILLER_176_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18234_ _02491_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__clkbuf_1
X_15446_ rbzero.wall_tracer.visualWallDist\[3\] _08475_ vssd1 vssd1 vccd1 vccd1 _08541_
+ sky130_fd_sc_hd__nand2_2
X_12658_ _05648_ _04657_ _05822_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__mux2_1
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18165_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__and2_1
X_11609_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__inv_2
XFILLER_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15377_ rbzero.wall_tracer.visualWallDist\[-11\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _08472_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12589_ _05764_ _05766_ _05767_ _05768_ net20 vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a32o_1
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _10136_ sky130_fd_sc_hd__or2_1
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _07438_ _07439_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__xnor2_1
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18096_ _02374_ _02375_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__nor2_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17047_ _10066_ _10067_ vssd1 vssd1 vccd1 vccd1 _10068_ sky130_fd_sc_hd__xor2_1
XFILLER_172_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03785_ _03785_ vssd1 vssd1 vccd1 vccd1 clknet_0__03785_ sky130_fd_sc_hd__clkbuf_16
X_14259_ _07367_ _07421_ _07428_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__nand3_1
XFILLER_131_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _08116_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17949_ _02235_ _02236_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__or2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20960_ clknet_leaf_64_i_clk _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ rbzero.pov.ss_buffer\[1\] _04052_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__nor2_2
X_20891_ clknet_leaf_44_i_clk _00480_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_4
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21512_ clknet_leaf_81_i_clk _01101_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21443_ net161 _01032_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21374_ clknet_leaf_24_i_clk _00963_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20313__177 clknet_1_0__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__inv_2
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20187_ _03384_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__buf_4
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19650__32 clknet_1_0__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11960_ rbzero.debug_overlay.facingX\[-5\] _05112_ _05064_ vssd1 vssd1 vccd1 vccd1
+ _05149_ sky130_fd_sc_hd__a21bo_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10911_ _04251_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _05078_ _05079_ _04638_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand3b_4
X_13630_ _06799_ _06800_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__xor2_1
X_10842_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__clkbuf_4
X_20563__23 clknet_1_0__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XFILLER_38_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ _06633_ _06696_ _06699_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__a21oi_4
X_10773_ rbzero.tex_g1\[16\] rbzero.tex_g1\[17\] _04177_ vssd1 vssd1 vccd1 vccd1 _04179_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15300_ rbzero.side_hot vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__inv_2
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _05661_ net8 vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__nor2_1
X_16280_ _09370_ _09371_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13492_ _06618_ _06576_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__nand2_1
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15231_ _08276_ _08314_ _08325_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__or3_1
X_12443_ _05263_ _05555_ _05557_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a31o_1
XFILLER_200_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ _08256_ rbzero.debug_overlay.playerX\[-4\] _08185_ vssd1 vssd1 vccd1 vccd1
+ _08257_ sky130_fd_sc_hd__mux2_1
X_12374_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _04931_ vssd1 vssd1 vccd1 vccd1 _05559_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ _07257_ _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__xnor2_2
XFILLER_176_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11325_ _04473_ _04513_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21a_1
X_19970_ _08220_ _03611_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nand2_1
X_15093_ rbzero.debug_overlay.playerX\[-8\] _08185_ vssd1 vssd1 vccd1 vccd1 _08188_
+ sky130_fd_sc_hd__nand2_1
XFILLER_158_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14044_ _07166_ _07197_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__and2b_2
X_18921_ _03042_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
X_11256_ gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__nand2_2
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11187_ rbzero.tex_b0\[12\] rbzero.tex_b0\[11\] _04395_ vssd1 vssd1 vccd1 vccd1 _04396_
+ sky130_fd_sc_hd__mux2_1
X_18852_ _03006_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
X_17803_ _01832_ _02029_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__and2_1
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18783_ _02970_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15995_ _08572_ _08613_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__nor2_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17734_ _02005_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__xnor2_1
X_14946_ _08065_ _08077_ _08078_ _08061_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__o211a_1
XFILLER_36_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _01828_ _01847_ _01845_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14877_ _08028_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16616_ _09575_ _09576_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__nor2_1
X_19404_ _03324_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
X_13828_ _06996_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__nand2_1
XFILLER_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17596_ _01885_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__nand2_1
XFILLER_165_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16547_ _09635_ _09636_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__and2b_1
X_19335_ rbzero.spi_registers.new_sky\[2\] rbzero.spi_registers.got_new_sky _03097_
+ _04409_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a31o_1
X_13759_ _06928_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nand2b_1
XFILLER_188_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19266_ rbzero.spi_registers.texadd3\[2\] _03242_ vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__or2_1
XFILLER_206_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16478_ _09561_ _09568_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__xnor2_2
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _02480_ vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__clkbuf_1
X_15429_ _08521_ _08523_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__xor2_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19197_ rbzero.spi_registers.new_texadd\[1\]\[22\] _03173_ _03203_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__o211a_1
XFILLER_129_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03806_ clknet_0__03806_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03806_
+ sky130_fd_sc_hd__clkbuf_16
X_18148_ _02419_ _02414_ _02417_ _02418_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__o211ai_2
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18079_ _02359_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__or2b_1
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20110_ rbzero.pov.ready_buffer\[6\] _03663_ _03709_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01236_ sky130_fd_sc_hd__o211a_1
X_21090_ clknet_leaf_97_i_clk _00679_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20041_ rbzero.debug_overlay.facingX\[-1\] _03663_ _03671_ _03669_ vssd1 vssd1 vccd1
+ vccd1 _01205_ sky130_fd_sc_hd__a211o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21992_ net138 _01581_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20943_ clknet_leaf_52_i_clk _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20874_ clknet_leaf_19_i_clk _00463_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_hot\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21426_ clknet_leaf_95_i_clk _01015_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21357_ clknet_leaf_21_i_clk _00946_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11110_ _04355_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12090_ _04656_ _04704_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__xnor2_1
X_21288_ clknet_leaf_6_i_clk _00877_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11041_ _04319_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__05993_ clknet_0__05993_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05993_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _07866_ _07958_ _07963_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__nand3_2
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _08039_ _08847_ _08274_ _08458_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__nor4_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ rbzero.wall_tracer.trackDistX\[6\] vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__inv_2
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14731_ _07899_ _07804_ _07827_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__mux2_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ rbzero.debug_overlay.vplaneY\[-4\] vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__buf_2
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17450_ _10308_ _10357_ _10355_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a21oi_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14662_ _07407_ _07832_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__xnor2_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11874_ _04824_ _05062_ _04424_ _03977_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__or4bb_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20476__324 clknet_1_1__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__inv_2
X_16401_ _08616_ _09489_ _09491_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__nor3_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _06771_ _06783_ _06754_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__or3_1
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10825_ rbzero.tex_g0\[56\] rbzero.tex_g0\[55\] _04203_ vssd1 vssd1 vccd1 vccd1 _04206_
+ sky130_fd_sc_hd__mux2_1
X_17381_ _10289_ _10312_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__or2b_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ _07760_ _07761_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__or2_1
XFILLER_164_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19120_ rbzero.spi_registers.new_texadd\[0\]\[12\] _03155_ _03160_ _03158_ vssd1
+ vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__o211a_1
XFILLER_198_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16332_ _08012_ _08023_ _08450_ _09188_ _08027_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__o41a_1
X_13544_ _06595_ _06697_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__nor2_1
XFILLER_185_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10756_ rbzero.tex_g1\[24\] rbzero.tex_g1\[25\] _04166_ vssd1 vssd1 vccd1 vccd1 _04170_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19051_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__buf_2
XFILLER_200_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16263_ _09344_ _09346_ _09342_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__a21boi_4
XFILLER_187_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13475_ _06582_ _06590_ _06598_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__o211a_1
X_10687_ _04133_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__clkbuf_1
X_18002_ _02287_ _02288_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15214_ rbzero.debug_overlay.playerY\[-2\] _08281_ vssd1 vssd1 vccd1 vccd1 _08309_
+ sky130_fd_sc_hd__xor2_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12426_ _05609_ _05610_ _04826_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__mux2_1
X_16194_ _09270_ _09286_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20567__3 clknet_1_1__leaf__03457_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
X_15145_ _08239_ rbzero.debug_overlay.playerX\[-5\] _08218_ vssd1 vssd1 vccd1 vccd1
+ _08240_ sky130_fd_sc_hd__mux2_1
XFILLER_154_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _05017_ _05506_ _05539_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a31o_1
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _04489_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and2b_1
X_15076_ rbzero.wall_tracer.stepDistY\[-11\] _08149_ _06262_ _08170_ vssd1 vssd1 vccd1
+ vccd1 _08171_ sky130_fd_sc_hd__o211ai_4
X_19953_ _06133_ _03604_ _03437_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a21o_1
X_12288_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _05009_ vssd1 vssd1 vccd1 vccd1 _05474_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14027_ _07166_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__xnor2_2
XFILLER_49_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18904_ rbzero.pov.spi_buffer\[59\] rbzero.pov.ready_buffer\[59\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
X_11239_ _04433_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__buf_4
X_19884_ _03554_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ _02997_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15978_ _09071_ _09072_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__and2b_1
X_18766_ _02929_ _02957_ _02958_ _02952_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__a211oi_1
XFILLER_209_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17717_ rbzero.wall_tracer.visualWallDist\[4\] _08421_ vssd1 vssd1 vccd1 vccd1 _02007_
+ sky130_fd_sc_hd__nand2_1
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ rbzero.wall_tracer.visualWallDist\[-1\] _08046_ vssd1 vssd1 vccd1 vccd1 _08067_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18697_ _02895_ _02896_ _02879_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__o21bai_1
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17648_ _01937_ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__nand2_1
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17579_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nor2_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19318_ rbzero.floor_leak\[1\] _03272_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__or2_1
XFILLER_182_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20590_ _03820_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19249_ rbzero.spi_registers.texadd2\[20\] _03207_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__or2_1
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21211_ clknet_leaf_2_i_clk _00800_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21142_ clknet_leaf_10_i_clk _00731_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21073_ clknet_leaf_81_i_clk _00662_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20024_ rbzero.debug_overlay.facingX\[-7\] _03658_ vssd1 vssd1 vccd1 vccd1 _03661_
+ sky130_fd_sc_hd__or2_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20425__278 clknet_1_0__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__inv_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21975_ net501 _01564_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20926_ clknet_leaf_55_i_clk _00515_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ clknet_leaf_58_i_clk _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ rbzero.tex_r0\[30\] rbzero.tex_r0\[29\] _04088_ vssd1 vssd1 vccd1 vccd1 _04093_
+ sky130_fd_sc_hd__mux2_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ _04776_ _04775_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__nand2_1
XFILLER_195_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20788_ _03110_ _03963_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and3_1
XFILLER_70_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _04055_ vssd1 vssd1 vccd1 vccd1 _04057_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ _06332_ _06345_ _06409_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__and3_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20319__183 clknet_1_1__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__inv_2
X_10472_ _04018_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12211_ rbzero.tex_g1\[1\] _04904_ _05182_ _04918_ vssd1 vssd1 vccd1 vccd1 _05398_
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21409_ clknet_leaf_24_i_clk _00998_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _06305_ _06307_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _05328_ _05329_ _04947_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__mux2_1
XFILLER_159_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12073_ _04903_ _05248_ _05252_ _04887_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a311o_1
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16950_ _09689_ _09971_ _09045_ vssd1 vssd1 vccd1 vccd1 _09972_ sky130_fd_sc_hd__a21o_1
XFILLER_173_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11024_ _04310_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
X_15901_ _08763_ _08995_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__xnor2_2
X_16881_ _09901_ _09902_ vssd1 vssd1 vccd1 vccd1 _09903_ sky130_fd_sc_hd__xor2_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15832_ _08434_ _08696_ _08913_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__o21bai_1
X_18620_ _02809_ _02813_ _02823_ _02824_ _08136_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a311oi_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _08837_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__xnor2_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _02758_ _02759_ _02760_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__o21ai_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12975_ _06142_ _06143_ _06149_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__and4bb_2
XFILLER_205_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _01785_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__xnor2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14714_ _06579_ _07808_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__nor2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _02705_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
X_11926_ _05082_ _05093_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__nor2_4
X_15694_ _08732_ _08733_ _08788_ _08735_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__a22o_1
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _01717_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14645_ _07815_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__clkinv_2
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11857_ _04696_ _04697_ _04701_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__nor3_2
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17364_ _10284_ _10285_ _10282_ _10283_ vssd1 vssd1 vccd1 vccd1 _10382_ sky130_fd_sc_hd__o2bb2a_1
X_10808_ net50 rbzero.tex_g0\[63\] _04121_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14576_ _07716_ _07742_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__nor2_1
XFILLER_207_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11788_ _04913_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__buf_6
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16315_ _09170_ _09293_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__nand2_1
X_19103_ rbzero.spi_registers.new_texadd\[0\]\[5\] _03141_ _03150_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00788_ sky130_fd_sc_hd__o211a_1
XFILLER_174_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13527_ _06595_ _06697_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__nand2_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17295_ _08399_ _08553_ _10313_ vssd1 vssd1 vccd1 vccd1 _10314_ sky130_fd_sc_hd__or3_1
X_10739_ rbzero.tex_g1\[32\] rbzero.tex_g1\[33\] _04155_ vssd1 vssd1 vccd1 vccd1 _04161_
+ sky130_fd_sc_hd__mux2_1
XFILLER_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19034_ rbzero.spi_registers.new_other\[0\] _03098_ _03108_ _03103_ vssd1 vssd1 vccd1
+ vccd1 _00761_ sky130_fd_sc_hd__o211a_1
X_16246_ _09086_ _09220_ _09219_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19678__57 clknet_1_1__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
X_13458_ _06474_ _06510_ _06512_ _06508_ _06590_ _06576_ vssd1 vssd1 vccd1 vccd1 _06629_
+ sky130_fd_sc_hd__mux4_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12409_ rbzero.tex_b1\[11\] rbzero.tex_b1\[10\] _05314_ vssd1 vssd1 vccd1 vccd1 _05594_
+ sky130_fd_sc_hd__mux2_1
X_16177_ _09169_ _09173_ _09269_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ _06512_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__inv_2
XFILLER_86_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20530__373 clknet_1_0__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__inv_2
XFILLER_115_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15128_ _08221_ _08222_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19936_ _04674_ _03591_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nand2_1
X_15059_ _08147_ _08153_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__or2_1
XFILLER_123_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19867_ rbzero.pov.spi_buffer\[70\] rbzero.pov.spi_buffer\[71\] _03467_ vssd1 vssd1
+ vccd1 vccd1 _03546_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18818_ _02988_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19798_ rbzero.pov.spi_buffer\[37\] rbzero.pov.spi_buffer\[38\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XFILLER_68_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18749_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__or2_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21760_ net286 _01349_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20711_ _03922_ _04437_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__mux2_1
XFILLER_52_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21691_ net217 _01280_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20642_ _03860_ _03864_ _03865_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__o211a_1
XFILLER_165_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20573_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__or2_1
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21125_ clknet_leaf_92_i_clk _00714_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21056_ clknet_leaf_99_i_clk _00645_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__05761_ clknet_0__05761_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05761_
+ sky130_fd_sc_hd__clkbuf_16
X_20007_ _03640_ _04667_ _04673_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__and3b_1
XFILLER_59_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12760_ _05890_ _05936_ _05937_ _05551_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__o22a_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ net484 _01547_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ rbzero.color_sky\[0\] rbzero.color_floor\[0\] _04825_ vssd1 vssd1 vccd1 vccd1
+ _04901_ sky130_fd_sc_hd__mux2_1
XFILLER_187_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20909_ clknet_leaf_36_i_clk _00498_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12691_ net53 _05843_ _05845_ net55 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a22o_1
XFILLER_199_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21889_ net415 _01478_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _07598_ _07600_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__nor2_1
X_11642_ _04810_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__inv_4
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _07045_ _07248_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__or2_1
XFILLER_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _04763_ sky130_fd_sc_hd__and2_1
XFILLER_122_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16100_ rbzero.wall_tracer.stepDistY\[6\] _08405_ vssd1 vssd1 vccd1 vccd1 _09194_
+ sky130_fd_sc_hd__nand2_1
Xinput18 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ _06480_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nor2_1
X_17080_ _10087_ _10100_ vssd1 vssd1 vccd1 vccd1 _10101_ sky130_fd_sc_hd__xnor2_1
X_10524_ _04045_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__clkbuf_1
Xinput29 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14292_ _07452_ _07457_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__or2b_1
XFILLER_182_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16031_ _09000_ _09100_ _09098_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__a21boi_2
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ _06324_ _06328_ _06410_ _06322_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__a31o_1
XFILLER_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10455_ _04009_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ _06336_ _06338_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12125_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _05002_ vssd1 vssd1 vccd1 vccd1 _05313_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17982_ _02262_ _02269_ rbzero.wall_tracer.trackDistX\[9\] _09879_ vssd1 vssd1 vccd1
+ vccd1 _00548_ sky130_fd_sc_hd__o2bb2a_1
X_19721_ rbzero.pov.spi_buffer\[0\] rbzero.pov.spi_buffer\[1\] _03468_ vssd1 vssd1
+ vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XFILLER_46_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16933_ _09557_ _09667_ _09673_ _09663_ vssd1 vssd1 vccd1 vccd1 _09955_ sky130_fd_sc_hd__a22o_1
X_12056_ rbzero.tex_r1\[62\] _05031_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__or2_1
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _04301_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16864_ _06104_ _09721_ vssd1 vssd1 vccd1 vccd1 _09887_ sky130_fd_sc_hd__nand2_1
XFILLER_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18603_ _05127_ rbzero.wall_tracer.rayAddendY\[1\] vssd1 vssd1 vccd1 vccd1 _02809_
+ sky130_fd_sc_hd__nand2_1
X_15815_ _08410_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__clkbuf_4
X_16795_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09825_ sky130_fd_sc_hd__or2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19583_ _03382_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__buf_4
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15746_ _08840_ _08786_ _08793_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__nand3_1
X_18534_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__nor2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _04674_ rbzero.map_rom.f2 rbzero.wall_tracer.mapX\[5\] _06133_ vssd1 vssd1
+ vccd1 vccd1 _06134_ sky130_fd_sc_hd__a22o_1
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ _05093_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nor2_1
X_15677_ _08720_ _08721_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__xnor2_1
X_18465_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _02598_
+ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12889_ _06064_ _06014_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__xnor2_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17416_ _10190_ _10318_ _10320_ _10321_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22oi_2
X_14628_ _07578_ _07627_ _07796_ _07798_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__a22o_1
X_18396_ _02624_ _02613_ _02625_ _08134_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a31o_1
XFILLER_159_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17347_ _10144_ _10365_ vssd1 vssd1 vccd1 vccd1 _10366_ sky130_fd_sc_hd__nand2_1
XFILLER_187_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14559_ _07692_ _07729_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _10290_ _10186_ _10295_ vssd1 vssd1 vccd1 vccd1 _10297_ sky130_fd_sc_hd__and3_1
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ _09319_ _09321_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__xor2_1
X_19017_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__buf_4
XFILLER_177_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19919_ rbzero.pov.ready_buffer\[66\] _03438_ _03558_ _03580_ vssd1 vssd1 vccd1 vccd1
+ _03581_ sky130_fd_sc_hd__a211o_1
XFILLER_25_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21812_ net338 _01401_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21743_ net269 _01332_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21674_ clknet_leaf_7_i_clk _01263_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20537__379 clknet_1_1__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__inv_2
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20625_ _03851_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20236__107 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__inv_2
XFILLER_165_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20556_ clknet_1_1__leaf__04634_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__buf_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19657__38 clknet_1_0__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
XFILLER_69_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21108_ clknet_leaf_89_i_clk _00697_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13930_ _07060_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21039_ clknet_leaf_78_i_clk _00628_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20282__149 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__inv_2
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ _07019_ _07020_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__or2_1
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15600_ _08662_ _08694_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__xor2_1
X_12812_ net41 _05263_ _05958_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__mux2_1
X_16580_ _08466_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__clkbuf_4
X_13792_ _06957_ _06958_ _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__nor3_1
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _08609_ _08615_ _08624_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__and3_1
X_12743_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__nor2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ rbzero.spi_registers.new_texadd\[2\]\[14\] rbzero.spi_registers.spi_buffer\[14\]
+ _02494_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_91_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15462_ _08235_ _08327_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__nor2_1
X_12674_ net49 _05845_ _05847_ _05852_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a22o_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17201_ _08581_ _09691_ _09973_ vssd1 vssd1 vccd1 vccd1 _10221_ sky130_fd_sc_hd__nor3b_4
XFILLER_31_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _07532_ _07583_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11625_ _04779_ _04785_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__nand2_1
X_18181_ _02447_ _02448_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__or2b_1
X_15393_ _08042_ _08428_ _08445_ _08484_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__a2bb2o_1
X_17132_ _09005_ _09491_ vssd1 vssd1 vccd1 vccd1 _10152_ sky130_fd_sc_hd__nor2_1
X_14344_ _07499_ _07514_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__nor2_1
XFILLER_155_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11556_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _04746_
+ sky130_fd_sc_hd__nand2_1
XFILLER_184_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ rbzero.tex_r1\[12\] rbzero.tex_r1\[13\] _04035_ vssd1 vssd1 vccd1 vccd1 _04037_
+ sky130_fd_sc_hd__mux2_1
X_17063_ _09406_ _09186_ vssd1 vssd1 vccd1 vccd1 _10084_ sky130_fd_sc_hd__nor2_1
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14275_ _07362_ _07445_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__nand2_1
XFILLER_144_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11487_ rbzero.debug_overlay.playerX\[3\] _04410_ _04578_ _04671_ _04676_ vssd1 vssd1
+ vccd1 vccd1 _04677_ sky130_fd_sc_hd__o221a_1
XFILLER_171_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16014_ rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerX\[-9\] _08138_
+ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__mux2_1
X_13226_ _06313_ _06394_ _06395_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__and3_1
X_10438_ _04000_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _06033_ _06030_ _06325_ _05995_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a311o_4
XFILLER_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _04436_ _04635_ _05056_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__o211ai_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _02251_ _02252_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__xor2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _06161_ _06263_ _04432_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__a21oi_2
XFILLER_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16916_ _09519_ _08620_ _09937_ vssd1 vssd1 vccd1 vccd1 _09938_ sky130_fd_sc_hd__or3_1
X_12039_ rbzero.tex_r1\[45\] _05199_ _05032_ _04890_ vssd1 vssd1 vccd1 vccd1 _05228_
+ sky130_fd_sc_hd__a31o_1
X_17896_ _02163_ _02165_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__or2_1
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19635_ rbzero.pov.spi_counter\[3\] rbzero.pov.spi_counter\[2\] _03442_ rbzero.pov.spi_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a31o_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16847_ _09871_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__clkbuf_1
X_20341__202 clknet_1_1__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__inv_2
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19566_ _03411_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16778_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ _09808_ _09809_ vssd1 vssd1 vccd1 vccd1 _09810_ sky130_fd_sc_hd__and4_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _09765_ _09773_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__or2b_1
XFILLER_179_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15729_ _08823_ _08774_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__nor2_1
XFILLER_55_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19497_ _03375_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_59_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18448_ _08135_ _02674_ _02675_ _09751_ rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a32o_1
XFILLER_22_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18379_ _02596_ rbzero.wall_tracer.rayAddendX\[2\] _02586_ vssd1 vssd1 vccd1 vccd1
+ _02611_ sky130_fd_sc_hd__o21bai_1
XFILLER_18_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21390_ clknet_leaf_10_i_clk _00979_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22011_ clknet_leaf_50_i_clk _01600_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03790_ clknet_0__03790_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03790_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21726_ net252 _01315_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21657_ clknet_leaf_44_i_clk _01246_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11410_ _04494_ _04495_ rbzero.texu_hot\[0\] vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a21o_1
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20608_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03838_
+ sky130_fd_sc_hd__nor2_1
X_12390_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _04931_ vssd1 vssd1 vccd1 vccd1 _05575_
+ sky130_fd_sc_hd__mux2_1
XFILLER_177_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21588_ clknet_leaf_92_i_clk _01177_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_193_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_85 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_85/HI o_rgb[12] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_96 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_96/HI zeros[3] sky130_fd_sc_hd__conb_1
XFILLER_153_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11341_ rbzero.spi_registers.texadd0\[17\] _04467_ _04532_ vssd1 vssd1 vccd1 vccd1
+ _04533_ sky130_fd_sc_hd__o21a_1
XFILLER_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ _07224_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11272_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__buf_4
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13011_ rbzero.wall_tracer.trackDistX\[-9\] vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__inv_2
XFILLER_134_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17750_ _02037_ _02038_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__and2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14962_ rbzero.wall_tracer.visualWallDist\[9\] _08047_ _08089_ _08085_ vssd1 vssd1
+ vccd1 vccd1 _00433_ sky130_fd_sc_hd__o211a_1
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ rbzero.traced_texa\[-5\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__a22o_1
X_13913_ _07075_ _07083_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__xor2_2
X_14893_ _08036_ _08038_ _08040_ _01633_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__o211a_1
XFILLER_130_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17681_ _01970_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__or2_1
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19420_ _02487_ rbzero.spi_registers.new_leak\[4\] _03329_ vssd1 vssd1 vccd1 vccd1
+ _03334_ sky130_fd_sc_hd__mux2_1
XFILLER_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ _06996_ _07006_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__xor2_1
X_16632_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerX\[-1\] _08138_
+ vssd1 vssd1 vccd1 vccd1 _09722_ sky130_fd_sc_hd__mux2_1
XFILLER_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19351_ rbzero.spi_registers.new_floor\[2\] _03289_ _03293_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00893_ sky130_fd_sc_hd__o211a_1
X_16563_ _09406_ _09176_ _09651_ _09652_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__o31a_1
XFILLER_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13775_ _06932_ _06945_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or2b_1
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10987_ rbzero.tex_b1\[42\] rbzero.tex_b1\[43\] _04281_ vssd1 vssd1 vccd1 vccd1 _04291_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18302_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__or2_1
XFILLER_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15514_ _08605_ _08606_ _08608_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__a21o_1
X_12726_ _05648_ _04657_ net28 vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__mux2_1
X_16494_ _09583_ _09584_ vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__xor2_1
X_19282_ rbzero.spi_registers.new_texadd\[3\]\[9\] _03240_ _03253_ _03252_ vssd1 vssd1
+ vccd1 vccd1 _00864_ sky130_fd_sc_hd__o211a_1
XFILLER_203_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15445_ _08538_ _08539_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__and2b_1
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18233_ rbzero.spi_registers.new_texadd\[2\]\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _02479_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
X_12657_ _05650_ _05651_ _05652_ _05653_ _05822_ net25 vssd1 vssd1 vccd1 vccd1 _05836_
+ sky130_fd_sc_hd__mux4_1
XFILLER_198_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11608_ _04751_ _04796_ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__or3_1
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15376_ _08042_ _08161_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__nor2_2
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18164_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nor2_1
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12588_ _05382_ _05470_ _05551_ _05632_ _05763_ net19 vssd1 vssd1 vccd1 vccd1 _05768_
+ sky130_fd_sc_hd__mux4_1
XFILLER_50_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17115_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _10135_ sky130_fd_sc_hd__nand2_1
X_14327_ _07479_ _07497_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__xnor2_1
X_11539_ _04723_ _04724_ _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__or3b_1
X_18095_ _02366_ _02368_ _02367_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a21boi_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17046_ _08535_ _09176_ vssd1 vssd1 vccd1 vccd1 _10067_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__03784_ _03784_ vssd1 vssd1 vccd1 vccd1 clknet_0__03784_ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14258_ _07367_ _07421_ _07428_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__a21o_1
XFILLER_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _06299_ _06300_ _06302_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__o21a_1
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _07160_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__or2_1
XFILLER_174_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _03083_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17948_ _02135_ _02145_ _02143_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a21oi_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17879_ _01878_ _02075_ _02073_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a21oi_2
XFILLER_54_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19618_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1
+ vccd1 _03439_ sky130_fd_sc_hd__nor2b_2
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20890_ clknet_leaf_45_i_clk _00479_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19549_ rbzero.spi_registers.new_texadd\[0\]\[16\] rbzero.spi_registers.spi_buffer\[16\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
XFILLER_206_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21511_ clknet_leaf_81_i_clk _01100_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_21442_ net160 _01031_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19714__89 clknet_1_0__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
XFILLER_148_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21373_ clknet_leaf_8_i_clk _00962_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20324_ clknet_1_1__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__buf_1
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20348__208 clknet_1_0__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__inv_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20186_ _03759_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10910_ rbzero.tex_g0\[16\] rbzero.tex_g0\[15\] _04248_ vssd1 vssd1 vccd1 vccd1 _04251_
+ sky130_fd_sc_hd__mux2_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11890_ _04415_ _04636_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__nand2_1
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _04053_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__buf_4
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13560_ _06687_ _06692_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__or2_1
X_10772_ _04178_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _05646_ _05057_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__or2_1
XFILLER_197_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21709_ net235 _01298_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _06619_ _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__or2_1
XFILLER_185_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15230_ _08318_ _08324_ _06263_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__mux2_4
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _05592_ _05626_ _05263_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a21oi_2
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15161_ _08254_ _08255_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__and2_1
X_12373_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _04931_ vssd1 vssd1 vccd1 vccd1 _05558_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ _07242_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__xor2_4
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ rbzero.spi_registers.texadd0\[13\] _04467_ _04515_ vssd1 vssd1 vccd1 vccd1
+ _04516_ sky130_fd_sc_hd__o21a_1
XFILLER_181_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15092_ _08185_ _08186_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__or2_1
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _07163_ _07198_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__nand2_2
X_18920_ rbzero.pov.spi_buffer\[67\] rbzero.pov.ready_buffer\[67\] _03033_ vssd1 vssd1
+ vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11255_ gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__or2_1
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20288__155 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__inv_2
XFILLER_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18851_ rbzero.pov.spi_buffer\[34\] rbzero.pov.ready_buffer\[34\] _03000_ vssd1 vssd1
+ vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
X_11186_ _04053_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__clkbuf_4
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17802_ _01842_ _02036_ _01839_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a21bo_1
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18782_ rbzero.pov.spi_buffer\[1\] rbzero.pov.ready_buffer\[1\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02970_ sky130_fd_sc_hd__mux2_1
X_15994_ _09073_ _09088_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__xnor2_2
XFILLER_209_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17733_ _02021_ _02022_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__nor2_1
XFILLER_48_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14945_ rbzero.wall_tracer.visualWallDist\[4\] _08046_ vssd1 vssd1 vccd1 vccd1 _08078_
+ sky130_fd_sc_hd__or2_1
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _01940_ _01954_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__xnor2_1
X_14876_ rbzero.wall_tracer.stepDistY\[8\] _08027_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08028_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19403_ _02487_ rbzero.spi_registers.new_floor\[4\] _03319_ vssd1 vssd1 vccd1 vccd1
+ _03324_ sky130_fd_sc_hd__mux2_1
X_16615_ _09661_ _09704_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13827_ _06995_ _06997_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__or2b_1
XFILLER_189_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17595_ _09519_ _09621_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__nor2_1
XFILLER_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19334_ rbzero.spi_registers.new_sky\[1\] _03280_ _03283_ _03278_ vssd1 vssd1 vccd1
+ vccd1 _00886_ sky130_fd_sc_hd__o211a_1
X_16546_ _09633_ _09634_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__nand2_1
X_13758_ _06888_ _06927_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__nand2_1
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12709_ _05882_ _05883_ _05885_ _05886_ net32 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a32o_1
XFILLER_206_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19265_ rbzero.spi_registers.new_texadd\[3\]\[1\] _03240_ _03244_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00856_ sky130_fd_sc_hd__o211a_1
X_20453__303 clknet_1_0__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__inv_2
X_16477_ _09562_ _09567_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__xor2_2
X_13689_ _06858_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ rbzero.spi_registers.new_texadd\[2\]\[0\] _02473_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02480_ sky130_fd_sc_hd__mux2_1
X_15428_ _08522_ _08374_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19196_ rbzero.spi_registers.texadd1\[22\] _03175_ vssd1 vssd1 vccd1 vccd1 _03203_
+ sky130_fd_sc_hd__or2_1
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03805_ clknet_0__03805_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03805_
+ sky130_fd_sc_hd__clkbuf_16
X_18147_ _02417_ _02418_ _02419_ _02414_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a211o_1
X_15359_ _08144_ _08452_ _08453_ _08168_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__a31o_2
XFILLER_172_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18078_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__nand2_1
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17029_ _09911_ _09919_ _09918_ vssd1 vssd1 vccd1 vccd1 _10050_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ rbzero.pov.ready_buffer\[41\] _03288_ _03665_ vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__and3_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21991_ net137 _01580_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ clknet_leaf_54_i_clk _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20873_ clknet_leaf_43_i_clk _00462_ vssd1 vssd1 vccd1 vccd1 reg_rgb\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21425_ clknet_leaf_94_i_clk _01014_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21356_ clknet_leaf_21_i_clk _00945_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21287_ clknet_leaf_3_i_clk _00876_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ rbzero.tex_b1\[17\] rbzero.tex_b1\[18\] _04314_ vssd1 vssd1 vccd1 vccd1 _04319_
+ sky130_fd_sc_hd__mux2_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ rbzero.spi_registers.new_texadd\[3\]\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__mux2_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ rbzero.wall_tracer.trackDistX\[7\] vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__inv_2
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ rbzero.debug_overlay.vplaneY\[-8\] _05117_ _05118_ rbzero.debug_overlay.vplaneY\[-7\]
+ _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a221o_1
XFILLER_85_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14730_ _07836_ _07841_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__xnor2_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _07402_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__xnor2_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11873_ _04415_ _04632_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nor2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20402__257 clknet_1_0__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__inv_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _09490_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ _06662_ _06667_ _06670_ _06611_ _06525_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__a32oi_4
X_10824_ _04205_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__clkbuf_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17380_ _10291_ _10294_ _10292_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a21bo_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _07753_ _07759_ _07762_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13543_ _06480_ _06474_ _06508_ _06482_ _06579_ _06589_ vssd1 vssd1 vccd1 vccd1 _06714_
+ sky130_fd_sc_hd__mux4_1
X_16331_ _08026_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__inv_2
X_10755_ _04169_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19050_ rbzero.spi_registers.got_new_mapd _03096_ vssd1 vssd1 vccd1 vccd1 _03119_
+ sky130_fd_sc_hd__nand2_2
X_16262_ rbzero.texu_hot\[2\] _08145_ _09354_ _08085_ vssd1 vssd1 vccd1 vccd1 _00468_
+ sky130_fd_sc_hd__o211a_1
X_13474_ _06521_ _06590_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__nand2_1
XFILLER_187_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ rbzero.tex_g1\[57\] rbzero.tex_g1\[58\] _04132_ vssd1 vssd1 vccd1 vccd1 _04133_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18001_ _09670_ _02012_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__nor2_1
X_15213_ _08307_ rbzero.debug_overlay.playerX\[-2\] _08218_ vssd1 vssd1 vccd1 vccd1
+ _08308_ sky130_fd_sc_hd__mux2_1
X_12425_ rbzero.tex_b1\[31\] rbzero.tex_b1\[30\] _04913_ vssd1 vssd1 vccd1 vccd1 _05610_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16193_ _09284_ _09285_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__and2_1
XFILLER_166_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15144_ rbzero.debug_overlay.playerX\[-5\] _08215_ vssd1 vssd1 vccd1 vccd1 _08239_
+ sky130_fd_sc_hd__xor2_1
X_12356_ _05029_ _05541_ _05043_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__o21ba_1
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ rbzero.texu_hot\[1\] _04492_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__a21o_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19952_ _06133_ _03605_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__nor2_1
X_15075_ _07867_ _08148_ _08169_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__a21o_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12287_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _05009_ vssd1 vssd1 vccd1 vccd1 _05473_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14026_ _07195_ _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__xnor2_2
X_18903_ _02966_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__buf_4
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11238_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__inv_4
XFILLER_106_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19883_ rbzero.pov.sclk_buffer\[1\] rbzero.pov.sclk_buffer\[0\] _03084_ vssd1 vssd1
+ vccd1 vccd1 _03554_ sky130_fd_sc_hd__mux2_1
XFILLER_150_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18834_ rbzero.pov.spi_buffer\[26\] rbzero.pov.ready_buffer\[26\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02997_ sky130_fd_sc_hd__mux2_1
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11169_ _04386_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18765_ rbzero.spi_registers.spi_counter\[2\] _02955_ rbzero.spi_registers.spi_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15977_ _09068_ _09070_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__nand2_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ _01897_ _01903_ _01902_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__o21ai_1
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14928_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.trackDistX\[-1\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__mux2_1
X_18696_ _02822_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02896_
+ sky130_fd_sc_hd__and2_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17647_ _01920_ _01921_ _01936_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__nand3_1
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _06600_ _07825_ _07866_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__o21ai_1
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17578_ _06169_ _09785_ _01869_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19317_ rbzero.spi_registers.new_leak\[0\] _03271_ _03273_ _03265_ vssd1 vssd1 vccd1
+ vccd1 _00879_ sky130_fd_sc_hd__o211a_1
X_16529_ _09365_ _09614_ _09492_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ rbzero.spi_registers.new_texadd\[2\]\[19\] _03221_ _03233_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__o211a_1
XFILLER_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19179_ rbzero.spi_registers.texadd1\[14\] _03189_ vssd1 vssd1 vccd1 vccd1 _03194_
+ sky130_fd_sc_hd__or2_1
XFILLER_157_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21210_ clknet_leaf_2_i_clk _00799_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21141_ clknet_leaf_7_i_clk _00730_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21072_ clknet_leaf_81_i_clk _00661_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20023_ rbzero.pov.ready_buffer\[34\] _03656_ _03660_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01198_ sky130_fd_sc_hd__o211a_1
XFILLER_59_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21974_ net500 _01563_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20925_ clknet_leaf_55_i_clk _00514_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20856_ clknet_leaf_58_i_clk _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20787_ gpout3.clk_div\[0\] gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__or2_1
XFILLER_23_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10540_ _04056_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10471_ rbzero.tex_r1\[29\] rbzero.tex_r1\[30\] _04013_ vssd1 vssd1 vccd1 vccd1 _04018_
+ sky130_fd_sc_hd__mux2_1
XFILLER_148_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ rbzero.tex_g1\[3\] _05305_ _05396_ _04947_ vssd1 vssd1 vccd1 vccd1 _05397_
+ sky130_fd_sc_hd__o211a_1
X_21408_ clknet_leaf_24_i_clk _00997_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13190_ _04427_ _06056_ _06360_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21o_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _05010_ vssd1 vssd1 vccd1 vccd1 _05329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21339_ clknet_leaf_9_i_clk _00928_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12072_ _05254_ _05256_ _05258_ _05260_ _04967_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__o221a_1
XFILLER_81_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11023_ rbzero.tex_b1\[25\] rbzero.tex_b1\[26\] _04303_ vssd1 vssd1 vccd1 vccd1 _04310_
+ sky130_fd_sc_hd__mux2_1
X_15900_ _08757_ _08811_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__nand2_1
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _09008_ _09490_ vssd1 vssd1 vccd1 vccd1 _09902_ sky130_fd_sc_hd__nor2_1
XFILLER_173_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _08921_ _08925_ _08923_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _02758_ _02759_ _02760_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__or3_1
XFILLER_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _08839_ _08855_ _08856_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__a21o_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _04720_ _04725_ rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _06150_
+ sky130_fd_sc_hd__a21o_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03808_ clknet_0__03808_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03808_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20326__188 clknet_1_1__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__inv_2
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _01786_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__xnor2_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _06613_ _07814_ _07882_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__o21bai_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _05111_ _05112_ _05113_ rbzero.debug_overlay.vplaneX\[-4\] _04652_ vssd1
+ vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a221o_1
X_18481_ _06088_ _02703_ _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XFILLER_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15693_ _08666_ _08734_ _08472_ _08457_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__or4_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17432_ _01719_ _01724_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__xor2_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11856_ _04900_ _04901_ _05018_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__o22a_1
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14644_ _07806_ _07814_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__or2_1
XFILLER_61_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _04196_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__clkbuf_1
X_17363_ _10307_ _10272_ vssd1 vssd1 vccd1 vccd1 _10381_ sky130_fd_sc_hd__or2b_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14575_ _07711_ _07743_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__nand2_1
X_11787_ _04958_ _04968_ _04976_ _04832_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a31o_1
XFILLER_202_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19102_ rbzero.spi_registers.texadd0\[5\] _03143_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__or2_1
XFILLER_186_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16314_ _08373_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__clkbuf_4
XFILLER_159_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10738_ _04160_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__clkbuf_1
X_13526_ _06585_ _06499_ _06501_ _06560_ _06554_ _06578_ vssd1 vssd1 vccd1 vccd1 _06697_
+ sky130_fd_sc_hd__mux4_1
X_17294_ _10289_ _10312_ vssd1 vssd1 vccd1 vccd1 _10313_ sky130_fd_sc_hd__xor2_1
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033_ rbzero.map_overlay.i_othery\[0\] _03101_ vssd1 vssd1 vccd1 vccd1 _03108_
+ sky130_fd_sc_hd__or2_1
X_16245_ _09239_ _09337_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13457_ _06495_ _06499_ _06501_ _06521_ _06590_ _06554_ vssd1 vssd1 vccd1 vccd1 _06628_
+ sky130_fd_sc_hd__mux4_1
X_10669_ rbzero.tex_r0\[2\] rbzero.tex_r0\[1\] _04121_ vssd1 vssd1 vccd1 vccd1 _04124_
+ sky130_fd_sc_hd__mux2_1
X_12408_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04978_ vssd1 vssd1 vccd1 vccd1 _05593_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16176_ _09174_ _09166_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__or2b_1
X_13388_ _06502_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__inv_2
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12339_ _05523_ _05524_ _04817_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__mux2_1
XFILLER_115_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ rbzero.debug_overlay.playerY\[-6\] _08202_ vssd1 vssd1 vccd1 vccd1 _08222_
+ sky130_fd_sc_hd__nand2_1
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19935_ rbzero.debug_overlay.playerX\[1\] _03559_ _03593_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01177_ sky130_fd_sc_hd__a211o_1
X_15058_ rbzero.wall_tracer.rayAddendY\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] _04463_
+ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__mux2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14009_ _07178_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__and2_1
X_19866_ _03545_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18817_ rbzero.pov.spi_buffer\[18\] rbzero.pov.ready_buffer\[18\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux2_1
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19797_ _03509_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18748_ rbzero.spi_registers.spi_counter\[4\] _02934_ vssd1 vssd1 vccd1 vccd1 _02944_
+ sky130_fd_sc_hd__or2_1
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18679_ _02821_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__and2_1
XFILLER_37_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20710_ _05050_ _03923_ _08045_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a21o_1
XFILLER_197_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21690_ net216 _01279_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20641_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03866_
+ sky130_fd_sc_hd__nand2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__05938_ clknet_0__05938_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05938_
+ sky130_fd_sc_hd__clkbuf_16
X_20572_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__nand2_1
XFILLER_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21124_ clknet_leaf_92_i_clk _00713_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21055_ clknet_leaf_95_i_clk _00644_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20006_ _03610_ _03643_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1
+ _03647_ sky130_fd_sc_hd__o21a_1
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21957_ net483 _01546_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__clkbuf_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ clknet_leaf_36_i_clk _00497_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ _05865_ _05868_ _05829_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__mux2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ net414 _01477_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ clknet_leaf_60_i_clk _00428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14360_ _07521_ _07519_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__xor2_2
X_11572_ _04759_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__nand2_1
XFILLER_156_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13311_ _06356_ _06481_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__xnor2_4
XFILLER_210_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10523_ rbzero.tex_r1\[4\] rbzero.tex_r1\[5\] _04035_ vssd1 vssd1 vccd1 vccd1 _04045_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_4
XFILLER_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14291_ _07414_ _07461_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__xnor2_1
X_20514__358 clknet_1_1__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__inv_2
XFILLER_196_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ _06330_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xor2_2
X_16030_ rbzero.texu_hot\[0\] _08145_ _09124_ _08085_ vssd1 vssd1 vccd1 vccd1 _00466_
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ rbzero.tex_r1\[37\] rbzero.tex_r1\[38\] _04002_ vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _04444_ _06341_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a21o_1
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _05310_ _05311_ _05191_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__mux2_1
X_17981_ _09872_ _02268_ _09879_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__o21a_1
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19720_ _03469_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
X_16932_ _09930_ _09953_ vssd1 vssd1 vccd1 vccd1 _09954_ sky130_fd_sc_hd__xnor2_1
X_12055_ _04903_ _05229_ _05233_ _04958_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a311o_1
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11006_ rbzero.tex_b1\[33\] rbzero.tex_b1\[34\] _04292_ vssd1 vssd1 vccd1 vccd1 _04301_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16863_ _09883_ _09884_ _09866_ vssd1 vssd1 vccd1 vccd1 _09886_ sky130_fd_sc_hd__a21o_1
XFILLER_81_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20408__263 clknet_1_1__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__inv_2
X_18602_ _02808_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15814_ _08898_ _08908_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__nand2_1
XFILLER_19_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19582_ _03419_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__clkbuf_1
X_16794_ _06187_ _09786_ _09824_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18533_ _02743_ _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__and2b_1
X_15745_ _08794_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__inv_2
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__inv_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ _02688_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nand2_1
X_11908_ _05083_ gpout0.hpos\[4\] _05075_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or3b_2
X_15676_ _08712_ _08766_ _08769_ _08770_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__nand2_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__xor2_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _07578_ _07627_ _07797_ _07579_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__a211oi_1
X_11839_ _05027_ rbzero.row_render.wall\[0\] _05026_ vssd1 vssd1 vccd1 vccd1 _05029_
+ sky130_fd_sc_hd__and3_1
X_18395_ _02624_ _02613_ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a21oi_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17346_ _10363_ _10364_ vssd1 vssd1 vccd1 vccd1 _10365_ sky130_fd_sc_hd__xor2_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14558_ _07423_ _07209_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__nor2_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13509_ _06589_ _06599_ _06679_ _06584_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__a22o_1
X_17277_ _10290_ _10186_ _10295_ vssd1 vssd1 vccd1 vccd1 _10296_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14489_ _07652_ _07653_ _07658_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__nand3_1
X_19016_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__buf_6
X_16228_ _09183_ _09202_ _09320_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _09131_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__buf_4
XFILLER_177_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19918_ _08307_ _03570_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nor2_1
XFILLER_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19849_ rbzero.pov.spi_buffer\[61\] rbzero.pov.spi_buffer\[62\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03537_ sky130_fd_sc_hd__mux2_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21811_ net337 _01400_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21742_ net268 _01331_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21673_ clknet_leaf_7_i_clk _01262_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20624_ _03844_ _03846_ _03845_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a21boi_1
XFILLER_149_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21107_ clknet_leaf_90_i_clk _00696_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21038_ clknet_leaf_79_i_clk _00627_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _07023_ _07029_ _07030_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12811_ _05952_ _05948_ _05983_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a31o_2
X_13791_ _06960_ _06961_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__xnor2_1
XFILLER_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15530_ _08609_ _08615_ _08624_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__a21oi_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _05899_ net28 vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__and2_1
XFILLER_128_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15461_ _08253_ _08328_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__nor2_1
X_12673_ _05711_ _05851_ net50 vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a21o_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _10096_ _10219_ vssd1 vssd1 vccd1 vccd1 _10220_ sky130_fd_sc_hd__xor2_1
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11624_ _04790_ _04806_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__or3_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _07253_ _07204_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__nor2_1
X_18180_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15392_ _08042_ _08428_ _08473_ _08445_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__or4b_1
X_20438__289 clknet_1_0__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__inv_2
X_17131_ _10031_ _10150_ vssd1 vssd1 vccd1 vccd1 _10151_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14343_ _07500_ _07512_ _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__a21oi_1
X_11555_ _04719_ _04742_ _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o21a_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ _04036_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17062_ _10077_ _10082_ vssd1 vssd1 vccd1 vccd1 _10083_ sky130_fd_sc_hd__xnor2_1
X_14274_ _07206_ _07444_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__nor2_1
X_11486_ _04672_ rbzero.debug_overlay.playerY\[3\] rbzero.debug_overlay.playerX\[2\]
+ _04421_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__o221a_1
XFILLER_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16013_ _08991_ _08993_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__xor2_4
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13225_ _06313_ _06394_ _06395_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10437_ rbzero.tex_r1\[45\] rbzero.tex_r1\[46\] _03991_ vssd1 vssd1 vccd1 vccd1 _04000_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ _05176_ _05295_ _05051_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__buf_6
X_17964_ _02158_ _02159_ _02161_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__o21a_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16915_ _09935_ _09936_ vssd1 vssd1 vccd1 vccd1 _09937_ sky130_fd_sc_hd__or2b_1
X_12038_ rbzero.tex_r1\[47\] _05002_ _05226_ _04922_ vssd1 vssd1 vccd1 vccd1 _05227_
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17895_ _02176_ _02183_ rbzero.wall_tracer.trackDistX\[8\] _09879_ vssd1 vssd1 vccd1
+ vccd1 _00547_ sky130_fd_sc_hd__o2bb2a_1
X_19634_ rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\] _03448_ vssd1 vssd1
+ vccd1 vccd1 _03451_ sky130_fd_sc_hd__and3_1
X_16846_ rbzero.wall_tracer.trackDistX\[-3\] _09870_ _09844_ vssd1 vssd1 vccd1 vccd1
+ _09871_ sky130_fd_sc_hd__mux2_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19565_ rbzero.spi_registers.new_texadd\[1\]\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
X_16777_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13989_ _07155_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ _09879_ _02730_ _02731_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a21oi_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15728_ _08246_ _08344_ _08719_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__nor3_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19496_ rbzero.spi_registers.new_mapd\[12\] rbzero.spi_registers.spi_buffer\[12\]
+ _03361_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _02672_ _02673_ _02668_ _02669_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a211o_1
X_15659_ _08727_ _08752_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__or2b_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18378_ rbzero.wall_tracer.rayAddendX\[2\] rbzero.wall_tracer.rayAddendX\[1\] _02596_
+ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ _10339_ _10347_ vssd1 vssd1 vccd1 vccd1 _10348_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22010_ clknet_leaf_37_i_clk _01599_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21725_ net251 _01314_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21656_ clknet_leaf_44_i_clk _01245_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20607_ rbzero.texV\[-6\] _03695_ _03819_ _03837_ vssd1 vssd1 vccd1 vccd1 _01605_
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21587_ clknet_leaf_92_i_clk _01176_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
Xtop_ew_algofoogle_75 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_75/HI o_rgb[0] sky130_fd_sc_hd__conb_1
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_86 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_86/HI o_rgb[13] sky130_fd_sc_hd__conb_1
XFILLER_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ rbzero.spi_registers.texadd1\[17\] _04461_ _04470_ _04531_ vssd1 vssd1 vccd1
+ vccd1 _04532_ sky130_fd_sc_hd__a211o_1
Xtop_ew_algofoogle_97 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_97/HI zeros[4] sky130_fd_sc_hd__conb_1
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ rbzero.side_hot vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__buf_2
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ rbzero.wall_tracer.trackDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__inv_2
XFILLER_165_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14961_ rbzero.wall_tracer.trackDistX\[9\] _08037_ _08035_ _08088_ vssd1 vssd1 vccd1
+ vccd1 _08089_ sky130_fd_sc_hd__a211o_1
XFILLER_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16700_ rbzero.traced_texa\[-6\] _09755_ _09756_ rbzero.wall_tracer.visualWallDist\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13912_ _07081_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__nor2_1
XFILLER_48_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17680_ _10383_ _01859_ _01858_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a21oi_4
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14892_ _04442_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__buf_4
XFILLER_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16631_ _09602_ _09720_ vssd1 vssd1 vccd1 vccd1 _09721_ sky130_fd_sc_hd__xnor2_4
XFILLER_78_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ _07009_ _07013_ _06973_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__and3b_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19350_ rbzero.color_floor\[2\] _03290_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or2_1
X_16562_ _08813_ _09176_ _09037_ _09406_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__o22ai_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ _04290_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13774_ _06940_ _06943_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o21bai_1
X_18301_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__and2_1
X_15513_ _08545_ _08607_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__nand2_1
XFILLER_16_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12725_ _05901_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or2_1
X_19281_ rbzero.spi_registers.texadd3\[9\] _03242_ vssd1 vssd1 vccd1 vccd1 _03253_
+ sky130_fd_sc_hd__or2_1
X_16493_ _09384_ _09456_ _09454_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18232_ _02490_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15444_ _08164_ _08165_ _08537_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__or3b_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12656_ _05829_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__inv_2
XFILLER_157_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18163_ _01759_ _02433_ _02364_ rbzero.wall_tracer.trackDistY\[4\] vssd1 vssd1 vccd1
+ vccd1 _00565_ sky130_fd_sc_hd__o2bb2a_1
X_11607_ rbzero.texV\[7\] _04754_ _04753_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a21boi_1
X_15375_ _08429_ _08440_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__or2_2
X_12587_ _05763_ _05297_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__nand2_1
XFILLER_8_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20371__229 clknet_1_0__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__inv_2
XFILLER_168_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17114_ _06202_ _09785_ _10134_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14326_ _07481_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__xor2_1
XFILLER_144_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ rbzero.map_overlay.i_mapdx\[0\] _04413_ _03972_ _04726_ _04727_ vssd1 vssd1
+ vccd1 vccd1 _04728_ sky130_fd_sc_hd__o221a_1
X_18094_ _02372_ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__or2b_1
XFILLER_102_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17045_ _09942_ _10065_ vssd1 vssd1 vccd1 vccd1 _10066_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03783_ _03783_ vssd1 vssd1 vccd1 vccd1 clknet_0__03783_ sky130_fd_sc_hd__clkbuf_16
X_14257_ _07375_ _07376_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__xnor2_1
X_11469_ _04446_ _04448_ _04647_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _06378_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__clkinv_4
XFILLER_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _07155_ _07159_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__and2_1
XFILLER_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13139_ _06291_ _06296_ _06305_ _06309_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ net44 rbzero.spi_registers.mosi_buffer\[0\] _09734_ vssd1 vssd1 vccd1 vccd1
+ _03083_ sky130_fd_sc_hd__mux2_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _02233_ _02234_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__or2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20265__134 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__inv_2
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17878_ _01992_ _02166_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__xnor2_1
X_16829_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09855_ sky130_fd_sc_hd__nand2_1
X_19617_ rbzero.pov.spi_done rbzero.pov.ready _03118_ _03438_ vssd1 vssd1 vccd1 vccd1
+ _01014_ sky130_fd_sc_hd__o211a_1
XFILLER_94_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19548_ _03402_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _03366_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21510_ clknet_leaf_81_i_clk _01099_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21441_ net159 _01030_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21372_ clknet_leaf_20_i_clk _00961_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_mapd
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20323_ clknet_1_1__leaf__04634_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__buf_1
XFILLER_134_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20185_ rbzero.spi_registers.new_texadd\[3\]\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_90_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ _04213_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ rbzero.tex_g1\[17\] rbzero.tex_g1\[18\] _04177_ vssd1 vssd1 vccd1 vccd1 _04178_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _05661_ _05640_ _05666_ _05691_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a31o_2
X_21708_ net234 _01297_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
X_13490_ _06576_ _06659_ _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__o21a_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ _04887_ _05600_ _05608_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a31o_1
X_21639_ clknet_leaf_85_i_clk _01228_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ rbzero.row_render.texu\[0\] _05186_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_
+ sky130_fd_sc_hd__a21o_1
X_15160_ rbzero.debug_overlay.playerX\[-5\] _08215_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_43_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_166_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ _04514_ _04456_ _04462_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a21oi_1
X_14111_ _07280_ _07281_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__and2_1
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15091_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14042_ _07164_ _07198_ _07201_ _07162_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__a22o_2
X_11254_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__buf_4
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_58_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18850_ _03005_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11185_ _04394_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17801_ _02088_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__and2_1
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18781_ _02969_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
X_15993_ _09086_ _09087_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__nor2_1
X_17732_ _02019_ _02020_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__and2_1
X_14944_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.trackDistX\[4\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__mux2_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17663_ _01952_ _01953_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__nor2_1
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14875_ _07891_ _08026_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__or2_1
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19402_ _03323_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
X_16614_ _09701_ _09703_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__xnor2_1
X_13826_ _06952_ _06994_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__or2_1
X_17594_ _01776_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19333_ rbzero.color_sky\[1\] _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__or2_1
X_16545_ _09633_ _09634_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__nor2_1
X_13757_ _06888_ _06927_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__nor2_1
X_10969_ rbzero.tex_b1\[51\] rbzero.tex_b1\[52\] _04281_ vssd1 vssd1 vccd1 vccd1 _04282_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12708_ _05382_ _05470_ _05551_ _05632_ _05881_ net31 vssd1 vssd1 vccd1 vccd1 _05886_
+ sky130_fd_sc_hd__mux4_1
X_19264_ rbzero.spi_registers.texadd3\[1\] _03242_ vssd1 vssd1 vccd1 vccd1 _03244_
+ sky130_fd_sc_hd__or2_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16476_ _08039_ _08338_ _09566_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__or3_2
X_13688_ _06718_ _06798_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__or2_1
X_18215_ _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__buf_4
X_15427_ _08375_ _08372_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__and2_1
X_12639_ _05793_ _05803_ _05790_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nand3_1
XFILLER_15_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19195_ rbzero.spi_registers.new_texadd\[1\]\[21\] _03173_ _03202_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__o211a_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03804_ clknet_0__03804_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03804_
+ sky130_fd_sc_hd__clkbuf_16
X_18146_ _02411_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__inv_2
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15358_ _04464_ _06034_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__or2_2
XFILLER_141_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14309_ _07446_ _07451_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__nand2_1
X_18077_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__nor2_1
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15289_ _08383_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17028_ _10041_ _10048_ vssd1 vssd1 vccd1 vccd1 _10049_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ rbzero.spi_registers.spi_buffer\[20\] rbzero.spi_registers.spi_buffer\[19\]
+ _03051_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21990_ net136 _01579_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20941_ clknet_leaf_56_i_clk _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20872_ clknet_leaf_43_i_clk _00461_ vssd1 vssd1 vccd1 vccd1 reg_rgb\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21424_ clknet_leaf_6_i_clk _01013_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21355_ clknet_leaf_20_i_clk _00944_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_107_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21286_ clknet_leaf_3_i_clk _00875_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20168_ _03750_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__clkbuf_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20099_ rbzero.debug_overlay.vplaneY\[-8\] _03685_ vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__or2_1
X_12990_ rbzero.wall_tracer.trackDistY\[9\] _06162_ rbzero.wall_tracer.trackDistY\[8\]
+ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__a22o_1
XFILLER_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _05129_ _05121_ _05122_ rbzero.debug_overlay.vplaneY\[-9\] vssd1 vssd1 vccd1
+ vccd1 _05130_ sky130_fd_sc_hd__a22o_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _07828_ _07829_ _07830_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__o21a_1
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11872_ _04637_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__or2_2
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06766_ _06781_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nand2_1
X_10823_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _04203_ vssd1 vssd1 vccd1 vccd1 _04205_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14591_ _07760_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__nand2_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16330_ _09195_ _09421_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__and2_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13542_ _06619_ _06535_ _06653_ _06712_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__a31o_1
X_10754_ rbzero.tex_g1\[25\] rbzero.tex_g1\[26\] _04166_ vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16261_ _08145_ _09353_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__nand2_1
X_10685_ _03979_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__clkbuf_4
X_13473_ _06642_ _06643_ _06570_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__mux2_1
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20294__160 clknet_1_0__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__inv_2
X_18000_ _09662_ _02012_ _02229_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__o31a_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15212_ rbzero.debug_overlay.playerX\[-2\] _08277_ vssd1 vssd1 vccd1 vccd1 _08307_
+ sky130_fd_sc_hd__xor2_1
X_12424_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _04913_ vssd1 vssd1 vccd1 vccd1 _05609_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16192_ _09275_ _09283_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__or2_1
XFILLER_173_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _08214_ _08236_ _08237_ vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__a21bo_1
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _05019_ _05371_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__nand3_1
XFILLER_127_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ _04496_ _04497_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__nor2_1
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19951_ _03603_ _03606_ _03103_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__o21a_1
X_15074_ _08144_ _08167_ _08168_ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__a21o_1
X_12286_ rbzero.color_sky\[4\] rbzero.color_floor\[4\] _04825_ vssd1 vssd1 vccd1 vccd1
+ _05472_ sky130_fd_sc_hd__mux2_1
XFILLER_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14025_ _07094_ _07141_ _07139_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__a21oi_1
X_18902_ _03032_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
X_11237_ _04431_ _03974_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nand2_4
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19882_ _03553_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11168_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04384_ vssd1 vssd1 vccd1 vccd1 _04386_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18833_ _02996_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18764_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__and4_1
X_15976_ _09068_ _09070_ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__nor2_1
X_11099_ _04349_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17715_ _02003_ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__xor2_1
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ _08035_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__buf_2
XFILLER_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18695_ _02822_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02895_
+ sky130_fd_sc_hd__nor2_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ _01920_ _01921_ _01936_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a21o_1
XFILLER_1_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14858_ _08013_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _06975_ _06978_ _06979_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__a21oi_1
X_17577_ _09822_ _01764_ _01765_ _09812_ _01868_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__o311a_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14789_ _07947_ _07948_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__o21ai_4
X_20377__235 clknet_1_1__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__inv_2
X_19316_ rbzero.floor_leak\[0\] _03272_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__or2_1
XFILLER_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16528_ _09614_ _09617_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19247_ rbzero.spi_registers.texadd2\[19\] _03222_ vssd1 vssd1 vccd1 vccd1 _03233_
+ sky130_fd_sc_hd__or2_1
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16459_ _09406_ _09176_ _09549_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__or3_1
X_19178_ rbzero.spi_registers.new_texadd\[1\]\[13\] _03188_ _03193_ _03184_ vssd1
+ vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__o211a_1
XFILLER_118_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18129_ _02341_ _02403_ _02404_ _02339_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__o31a_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21140_ clknet_leaf_8_i_clk _00729_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21071_ clknet_leaf_81_i_clk _00660_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20022_ rbzero.debug_overlay.facingX\[-8\] _03658_ vssd1 vssd1 vccd1 vccd1 _03660_
+ sky130_fd_sc_hd__or2_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21973_ net499 _01562_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ clknet_leaf_56_i_clk _00513_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20855_ clknet_leaf_58_i_clk _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20786_ gpout3.clk_div\[0\] gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__nand2_1
XFILLER_167_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10470_ _04017_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21407_ clknet_leaf_24_i_clk _00996_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _04964_ vssd1 vssd1 vccd1 vccd1 _05328_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21338_ clknet_leaf_9_i_clk _00927_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ rbzero.tex_r1\[48\] _04982_ _04910_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_
+ sky130_fd_sc_hd__a31o_1
XFILLER_155_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21269_ clknet_leaf_28_i_clk _00858_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11022_ _04309_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _08923_ _08924_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__nor2_1
XFILLER_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _08841_ _08842_ _08854_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__and3_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12973_ _04721_ _06113_ _06145_ _06146_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__o221a_1
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03807_ clknet_0__03807_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03807_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _01790_ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__xor2_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14712_ _06579_ _07819_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__nor2_1
XFILLER_205_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _05089_ _05094_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nor2_4
X_18480_ _06161_ _06258_ _06264_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__o21a_2
X_15692_ _08235_ _08440_ _08736_ _08735_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__or4b_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17431_ _01722_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__xor2_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14643_ _07745_ _07788_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__xnor2_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _04900_ _05044_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__nand2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10806_ rbzero.tex_g1\[0\] rbzero.tex_g1\[1\] _04188_ vssd1 vssd1 vccd1 vccd1 _04196_
+ sky130_fd_sc_hd__mux2_1
X_17362_ _10377_ _10378_ _10261_ _10264_ vssd1 vssd1 vccd1 vccd1 _10380_ sky130_fd_sc_hd__a211oi_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14574_ _07714_ _07744_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__xor2_1
X_11786_ _04941_ _04971_ _04975_ _04902_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a211o_1
X_19101_ rbzero.spi_registers.new_texadd\[0\]\[4\] _03141_ _03149_ _03145_ vssd1 vssd1
+ vccd1 vccd1 _00787_ sky130_fd_sc_hd__o211a_1
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16313_ _09385_ _09404_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13525_ _06669_ _06694_ _06695_ _06651_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__o22a_1
X_10737_ rbzero.tex_g1\[33\] rbzero.tex_g1\[34\] _04155_ vssd1 vssd1 vccd1 vccd1 _04160_
+ sky130_fd_sc_hd__mux2_1
X_17293_ rbzero.wall_tracer.visualWallDist\[1\] _08475_ _08445_ vssd1 vssd1 vccd1
+ vccd1 _10312_ sky130_fd_sc_hd__and3_1
XFILLER_186_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ rbzero.spi_registers.new_other\[10\] _03098_ _03107_ _03103_ vssd1 vssd1
+ vccd1 vccd1 _00760_ sky130_fd_sc_hd__o211a_1
X_16244_ _09335_ _09336_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__nor2_1
X_13456_ _06619_ _06626_ _06602_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__o21ai_1
X_10668_ _04123_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _05565_ _05574_ _05582_ _05591_ _04810_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a221o_1
X_16175_ _09150_ _09160_ _09158_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__a21o_1
X_10599_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _04077_ vssd1 vssd1 vccd1 vccd1 _04087_
+ sky130_fd_sc_hd__mux2_1
X_13387_ _06493_ _06557_ _06530_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__or3b_2
XFILLER_86_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15126_ rbzero.debug_overlay.playerY\[-6\] _08202_ vssd1 vssd1 vccd1 vccd1 _08221_
+ sky130_fd_sc_hd__or2_1
XFILLER_99_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12338_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _04907_ vssd1 vssd1 vccd1 vccd1 _05524_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__clkbuf_4
X_19934_ rbzero.pov.ready_buffer\[69\] _03586_ _03591_ _03592_ _03569_ vssd1 vssd1
+ vccd1 vccd1 _03593_ sky130_fd_sc_hd__o221a_1
X_12269_ _04832_ _05437_ _05455_ net42 vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a31o_1
XFILLER_130_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14008_ _06540_ _06942_ _07177_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__o21ai_1
X_19865_ rbzero.pov.spi_buffer\[69\] rbzero.pov.spi_buffer\[70\] _03467_ vssd1 vssd1
+ vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
XFILLER_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03465_ _03465_ vssd1 vssd1 vccd1 vccd1 clknet_0__03465_ sky130_fd_sc_hd__clkbuf_16
X_18816_ _02987_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19796_ rbzero.pov.spi_buffer\[36\] rbzero.pov.spi_buffer\[37\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _08461_ _09053_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__nor2_1
X_18747_ rbzero.spi_registers.spi_counter\[0\] _02935_ _02941_ _02942_ rbzero.spi_registers.spi_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a32o_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18678_ _02821_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _02879_
+ sky130_fd_sc_hd__nor2_1
XFILLER_52_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17629_ _01831_ _01836_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__nand2_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20220__93 clknet_1_1__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
X_20640_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03865_
+ sky130_fd_sc_hd__or2_1
XFILLER_51_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20571_ gpout5.clk_div\[0\] net63 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__nor2_1
XFILLER_191_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20431__284 clknet_1_1__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__inv_2
XFILLER_132_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ clknet_leaf_91_i_clk _00712_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21054_ clknet_leaf_95_i_clk _00643_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20005_ rbzero.debug_overlay.playerY\[3\] _03611_ _03646_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01194_ sky130_fd_sc_hd__a211o_1
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21956_ net482 _01545_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ clknet_leaf_36_i_clk _00496_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_188_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ net413 _01476_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11640_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__buf_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20838_ clknet_leaf_65_i_clk _00427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _04757_ _04758_ rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a21o_1
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20769_ _02746_ _02751_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__and2b_1
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _06415_ _06392_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__nand2_2
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ _04044_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14290_ _07415_ _07441_ _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__o21a_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10453_ _04008_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__clkbuf_1
X_13241_ _06332_ _06345_ _06409_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__a31o_1
XFILLER_171_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13172_ _06327_ _06039_ _06040_ _06342_ _06323_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__o311a_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _04932_ vssd1 vssd1 vccd1 vccd1 _05311_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19683__62 clknet_1_1__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
X_17980_ _02265_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__xnor2_1
XFILLER_123_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16931_ _09932_ _09952_ vssd1 vssd1 vccd1 vccd1 _09953_ sky130_fd_sc_hd__xor2_1
X_12054_ _05235_ _05238_ _05240_ _05242_ _04967_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__o221a_1
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11005_ _04300_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16862_ _09883_ _09884_ vssd1 vssd1 vccd1 vccd1 _09885_ sky130_fd_sc_hd__nor2_1
XFILLER_93_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15813_ _08896_ _08897_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__or2_1
X_18601_ rbzero.wall_tracer.rayAddendY\[0\] _02807_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02808_ sky130_fd_sc_hd__mux2_1
X_19581_ rbzero.spi_registers.new_texadd\[1\]\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__mux2_1
X_16793_ _06105_ _09820_ _09821_ _09812_ _09823_ vssd1 vssd1 vccd1 vccd1 _09824_ sky130_fd_sc_hd__o311a_1
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18532_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__nand2_1
X_15744_ _08826_ _08838_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__xnor2_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12956_ rbzero.debug_overlay.playerY\[2\] _06086_ rbzero.map_rom.a6 _04667_ _06131_
+ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a221o_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _02598_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _02689_
+ sky130_fd_sc_hd__nand2_1
X_11907_ _05085_ _05093_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nor2_1
X_15675_ _08228_ _08298_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__nor2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12887_ _06013_ _06016_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__xor2_2
XFILLER_209_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _09397_ _09186_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__nor2_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14626_ _07577_ _07578_ _07627_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__nor3_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ rbzero.row_render.wall\[0\] rbzero.row_render.wall\[1\] _05023_ _05026_ _05027_
+ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a41o_1
X_18394_ _02596_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _02625_
+ sky130_fd_sc_hd__xor2_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17345_ _10146_ _10238_ _10236_ vssd1 vssd1 vccd1 vccd1 _10364_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14557_ _07417_ _07361_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__nor2_1
X_11769_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _04914_ vssd1 vssd1 vccd1 vccd1 _04959_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13508_ _06582_ _06504_ _06578_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__mux2_1
X_17276_ _10293_ _10294_ vssd1 vssd1 vccd1 vccd1 _10295_ sky130_fd_sc_hd__xor2_1
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14488_ _07652_ _07653_ _07658_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__a21o_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19015_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__buf_6
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16227_ _09197_ _09198_ _09201_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__and3_1
XFILLER_146_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ _06569_ _06538_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__nand2_1
XFILLER_173_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20489__336 clknet_1_1__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__inv_2
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _08304_ _09131_ _09250_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__or3_1
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _08202_ _08203_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__and2_1
XFILLER_177_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16089_ _09181_ _09182_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__nor2_1
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19917_ rbzero.debug_overlay.playerX\[-3\] _03569_ _03578_ _03579_ vssd1 vssd1 vccd1
+ vccd1 _01173_ sky130_fd_sc_hd__o211a_1
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19848_ _03536_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ rbzero.pov.spi_buffer\[28\] rbzero.pov.spi_buffer\[29\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03500_ sky130_fd_sc_hd__mux2_1
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21810_ net336 _01399_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21741_ net267 _01330_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21672_ clknet_leaf_26_i_clk _01261_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20623_ _03849_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__and2b_1
XFILLER_164_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21106_ clknet_leaf_70_i_clk _00695_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21037_ clknet_leaf_80_i_clk _00626_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _05946_ _05958_ _05985_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a31o_2
XFILLER_90_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ _06949_ _06953_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__and2_1
XFILLER_90_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _05711_ _05911_ _05917_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a31o_1
XFILLER_16_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21939_ net465 _01528_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _08552_ _08554_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__and2_1
XFILLER_31_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ net27 net26 vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__nor2_1
XFILLER_31_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _07534_ _07581_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__nand2_1
X_11623_ _04789_ _04778_ _04786_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__nor3_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _08470_ _08485_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__xor2_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17130_ _09525_ _09242_ vssd1 vssd1 vccd1 vccd1 _10150_ sky130_fd_sc_hd__nor2_1
XFILLER_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14342_ _07503_ _07511_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__and2b_1
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _04683_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__nor2_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10505_ rbzero.tex_r1\[13\] rbzero.tex_r1\[14\] _04035_ vssd1 vssd1 vccd1 vccd1 _04036_
+ sky130_fd_sc_hd__mux2_1
X_17061_ _09195_ _09421_ _08889_ vssd1 vssd1 vccd1 vccd1 _10082_ sky130_fd_sc_hd__a21oi_2
XFILLER_155_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14273_ _07443_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ gpout0.vpos\[7\] _04673_ _04674_ _04411_ vssd1 vssd1 vccd1 vccd1 _04675_
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _09105_ _09106_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__or2_1
X_13224_ _06286_ _06285_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__nand2_1
X_10436_ _03999_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13155_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__inv_2
XFILLER_100_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _04650_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__nor2_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17963_ _02245_ _02250_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__xor2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__buf_8
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16914_ _09933_ _09934_ vssd1 vssd1 vccd1 vccd1 _09936_ sky130_fd_sc_hd__nand2_1
X_12037_ rbzero.tex_r1\[46\] _05031_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__or2_1
XFILLER_78_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17894_ _02181_ _02182_ _09785_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19633_ rbzero.pov.spi_counter\[3\] _03448_ _03450_ _03446_ vssd1 vssd1 vccd1 vccd1
+ _01018_ sky130_fd_sc_hd__o211a_1
X_16845_ _09865_ _09867_ _09869_ vssd1 vssd1 vccd1 vccd1 _09870_ sky130_fd_sc_hd__o21ai_1
XFILLER_92_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16776_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09808_ sky130_fd_sc_hd__or2_1
X_19564_ _03410_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _07156_ _07158_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nor2_1
XFILLER_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15727_ _08287_ _08358_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__or2_1
X_18515_ rbzero.map_rom.f2 _09879_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__nor2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _04671_ _06113_ rbzero.wall_tracer.mapY\[5\] _06114_ vssd1 vssd1 vccd1 vccd1
+ _06115_ sky130_fd_sc_hd__a22o_1
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _03374_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15658_ _08727_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__xnor2_1
X_18446_ _02668_ _02669_ _02672_ _02673_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o211ai_2
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14609_ _07767_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18377_ _02596_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02609_
+ sky130_fd_sc_hd__nor2_1
X_15589_ _08681_ _08682_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__xor2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17328_ _10345_ _10346_ vssd1 vssd1 vccd1 vccd1 _10347_ sky130_fd_sc_hd__xor2_1
XFILLER_187_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17259_ _10150_ _10275_ _10277_ vssd1 vssd1 vccd1 vccd1 _10278_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19662__43 clknet_1_1__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
XFILLER_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20543__385 clknet_1_0__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__inv_2
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20242__113 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__inv_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ net250 _01313_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21655_ clknet_leaf_44_i_clk _01244_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_123_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20606_ _03835_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21586_ clknet_leaf_91_i_clk _01175_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_193_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_76 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_76/HI o_rgb[1] sky130_fd_sc_hd__conb_1
XFILLER_165_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_87 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_87/HI o_rgb[16] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_98 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_98/HI zeros[5] sky130_fd_sc_hd__conb_1
XFILLER_166_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20468_ clknet_1_1__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__buf_1
X_11270_ rbzero.spi_registers.texadd3\[13\] _04457_ _04461_ rbzero.spi_registers.texadd1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a22o_1
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14960_ _06215_ _06216_ rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1 vccd1
+ _08088_ sky130_fd_sc_hd__nor3b_1
X_22069_ clknet_leaf_40_i_clk _01658_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13911_ _07076_ _07077_ _07080_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__and3_1
XFILLER_48_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14891_ _08039_ _08035_ vssd1 vssd1 vccd1 vccd1 _08040_ sky130_fd_sc_hd__nand2_1
XFILLER_130_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16630_ _09587_ _09719_ vssd1 vssd1 vccd1 vccd1 _09720_ sky130_fd_sc_hd__xor2_4
X_13842_ _06963_ _07008_ _07005_ _07007_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__o211ai_1
XFILLER_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16561_ _08813_ _09037_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__or2_1
X_13773_ _06933_ _06934_ _06939_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__and3_1
X_10985_ rbzero.tex_b1\[43\] rbzero.tex_b1\[44\] _04281_ vssd1 vssd1 vccd1 vccd1 _04290_
+ sky130_fd_sc_hd__mux2_1
X_15512_ _08543_ _08544_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__or2_1
X_18300_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__nor2_1
X_12724_ gpout0.vpos\[0\] _05651_ _05652_ _05653_ net28 net31 vssd1 vssd1 vccd1 vccd1
+ _05902_ sky130_fd_sc_hd__mux4_1
X_19280_ rbzero.spi_registers.new_texadd\[3\]\[8\] _03240_ _03251_ _03252_ vssd1 vssd1
+ vccd1 vccd1 _00863_ sky130_fd_sc_hd__o211a_1
X_16492_ _09514_ _09582_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18231_ rbzero.spi_registers.new_texadd\[2\]\[5\] _02489_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_188_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15443_ _08164_ _08165_ _08537_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__o21ba_1
X_12655_ _04687_ _05644_ _05645_ _04642_ _05822_ _05829_ vssd1 vssd1 vccd1 vccd1 _05834_
+ sky130_fd_sc_hd__mux4_1
XFILLER_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18162_ _02341_ _02431_ _02432_ _02339_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__o31a_1
X_11606_ _04749_ _04750_ rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15374_ _08448_ _08468_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__xnor2_2
XFILLER_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12586_ _05765_ net20 vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nor2_1
X_17113_ _09782_ _10127_ _10133_ vssd1 vssd1 vccd1 vccd1 _10134_ sky130_fd_sc_hd__and3_1
XFILLER_8_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14325_ _07488_ _07494_ _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__o21a_1
XFILLER_102_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11537_ rbzero.map_overlay.i_mapdx\[3\] _04418_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__xnor2_1
X_18093_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__nand2_1
XFILLER_184_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17044_ _09044_ _09046_ _08813_ vssd1 vssd1 vccd1 vccd1 _10065_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__03782_ _03782_ vssd1 vssd1 vccd1 vccd1 clknet_0__03782_ sky130_fd_sc_hd__clkbuf_16
X_14256_ _07421_ _07422_ _07425_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a31o_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ _04657_ _04651_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nand2_1
XFILLER_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13207_ rbzero.wall_tracer.rcp_sel\[0\] _06366_ _06368_ _06373_ _06377_ vssd1 vssd1
+ vccd1 vccd1 _06378_ sky130_fd_sc_hd__a2111oi_4
XFILLER_171_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10419_ _03990_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14187_ _07343_ _07354_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xnor2_1
X_11399_ _04454_ _04510_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nand2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13138_ _06291_ _06307_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__and3b_1
XFILLER_140_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _03082_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__clkbuf_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _02226_ _02232_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__nor2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ rbzero.map_overlay.i_othery\[1\] _06089_ _06244_ vssd1 vssd1 vccd1 vccd1
+ _06245_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17877_ _02163_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__xor2_1
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19616_ _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__clkbuf_4
X_16828_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09854_ sky130_fd_sc_hd__or2_1
XFILLER_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19547_ rbzero.spi_registers.new_texadd\[0\]\[15\] rbzero.spi_registers.spi_buffer\[15\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__mux2_1
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16759_ rbzero.wall_tracer.mapX\[8\] _09786_ _09784_ _09794_ vssd1 vssd1 vccd1 vccd1
+ _00525_ sky130_fd_sc_hd__a22o_1
XFILLER_111_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19478_ rbzero.spi_registers.new_mapd\[3\] _02485_ _03362_ vssd1 vssd1 vccd1 vccd1
+ _03366_ sky130_fd_sc_hd__mux2_1
XFILLER_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18429_ _02644_ _02647_ _02645_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__o21bai_1
XFILLER_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21440_ net158 _01029_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21371_ clknet_leaf_12_i_clk _00960_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20184_ _03758_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _04143_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__clkbuf_4
XFILLER_197_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21707_ net233 _01296_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12440_ _04823_ _05616_ _05624_ _04832_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a31o_1
X_21638_ clknet_leaf_85_i_clk _01227_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12371_ rbzero.row_render.texu\[0\] _05186_ _05042_ vssd1 vssd1 vccd1 vccd1 _05556_
+ sky130_fd_sc_hd__o21ai_1
X_21569_ clknet_leaf_96_i_clk _01158_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14110_ _07236_ _07258_ _07279_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__or3_1
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11322_ rbzero.spi_registers.texadd2\[13\] vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__inv_2
XFILLER_154_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15090_ _06335_ _08182_ _08184_ _06426_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__a31o_2
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14041_ _07161_ _07202_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__or2_2
XFILLER_107_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11253_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__inv_2
XFILLER_10_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11184_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _04384_ vssd1 vssd1 vccd1 vccd1 _04394_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20249__119 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__inv_2
X_17800_ _02025_ _02086_ _02087_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nand3_1
X_15992_ _08568_ _09074_ _09085_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__and3_1
X_18780_ rbzero.pov.spi_buffer\[0\] rbzero.pov.ready_buffer\[0\] _02968_ vssd1 vssd1
+ vccd1 vccd1 _02969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17731_ _02019_ _02020_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__nor2_1
X_14943_ _08065_ _08075_ _08076_ _08061_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__o211a_1
XFILLER_76_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17662_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__and2_1
XFILLER_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14874_ _06568_ _07988_ _08025_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__o21a_1
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19401_ _02485_ rbzero.spi_registers.new_floor\[3\] _03319_ vssd1 vssd1 vccd1 vccd1
+ _03323_ sky130_fd_sc_hd__mux2_1
X_16613_ _09554_ _09574_ _09702_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__a21o_1
X_13825_ _06952_ _06994_ _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__or3b_1
XFILLER_63_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17593_ _10059_ _09243_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__nor2_1
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20554__15 clknet_1_0__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16544_ _09497_ _09505_ _09503_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19332_ rbzero.spi_registers.got_new_sky _03096_ vssd1 vssd1 vccd1 vccd1 _03282_
+ sky130_fd_sc_hd__and2_1
X_13756_ _06924_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__and2b_1
X_10968_ _04143_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12707_ _05884_ net32 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__nor2_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19263_ rbzero.spi_registers.new_texadd\[3\]\[0\] _03240_ _03243_ _03237_ vssd1 vssd1
+ vccd1 vccd1 _00855_ sky130_fd_sc_hd__o211a_1
X_16475_ _08148_ _09564_ _09565_ _08454_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__a31o_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13687_ _06722_ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__nor2_1
XFILLER_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _04237_ vssd1 vssd1 vccd1 vccd1 _04245_
+ sky130_fd_sc_hd__mux2_1
XFILLER_148_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15426_ _08509_ _08511_ _08508_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__a21bo_1
X_18214_ _02474_ _02477_ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1
+ _02478_ sky130_fd_sc_hd__nor3b_4
X_12638_ _05779_ _05788_ _05813_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__or4b_2
X_19194_ rbzero.spi_registers.texadd1\[21\] _03175_ vssd1 vssd1 vccd1 vccd1 _03202_
+ sky130_fd_sc_hd__or2_1
XFILLER_54_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03803_ clknet_0__03803_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03803_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18145_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__or2_1
X_15357_ _04464_ _06426_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__nand2_1
XFILLER_145_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12569_ _04446_ _05715_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__nand2_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14308_ _07446_ _07478_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__nand2_1
X_18076_ _09830_ _02358_ _02340_ rbzero.wall_tracer.trackDistY\[-8\] vssd1 vssd1 vccd1
+ vccd1 _00553_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15288_ rbzero.wall_tracer.stepDistX\[-2\] _08162_ _08382_ vssd1 vssd1 vccd1 vccd1
+ _08383_ sky130_fd_sc_hd__a21boi_2
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17027_ _10042_ _10047_ vssd1 vssd1 vccd1 vccd1 _10048_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14239_ _07407_ _07408_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__and2_1
XFILLER_113_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _03073_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20460__309 clknet_1_1__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__inv_2
X_20227__99 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__inv_2
X_17929_ rbzero.wall_tracer.visualWallDist\[8\] _10183_ _01699_ rbzero.wall_tracer.visualWallDist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
XFILLER_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20940_ clknet_leaf_56_i_clk _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20871_ clknet_leaf_43_i_clk _00460_ vssd1 vssd1 vccd1 vccd1 reg_rgb\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20354__214 clknet_1_1__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__inv_2
XFILLER_148_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21423_ clknet_leaf_25_i_clk _01012_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21354_ clknet_leaf_20_i_clk _00943_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21285_ clknet_leaf_3_i_clk _00874_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20167_ _03732_ _03748_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__and3_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ rbzero.pov.ready_buffer\[0\] _03684_ _03702_ _03703_ vssd1 vssd1 vccd1 vccd1
+ _01230_ sky130_fd_sc_hd__o211a_1
XFILLER_188_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11871_ _04412_ _04636_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__nor2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13610_ _06779_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__nor2_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _04204_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _07752_ _07759_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__xnor2_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _06641_ _06695_ _06636_ _06577_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__a221o_1
X_10753_ _04168_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16260_ _09121_ _09352_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13472_ _06474_ _06510_ _06603_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__mux2_1
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _04131_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _08172_ _08305_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__nand2_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _04953_ _05603_ _05607_ _04902_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a211o_1
X_16191_ _09275_ _09283_ vssd1 vssd1 vccd1 vccd1 _09284_ sky130_fd_sc_hd__nand2_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15142_ _08178_ _08213_ _08195_ _08201_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__or4_1
XFILLER_154_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12354_ _05038_ _05372_ _05177_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a21o_1
XFILLER_153_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11305_ rbzero.texu_hot\[1\] _04492_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19950_ rbzero.pov.ready_buffer\[72\] _03586_ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_
+ sky130_fd_sc_hd__o21a_1
X_15073_ _04436_ rbzero.trace_state\[0\] _06259_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__and3_2
XFILLER_153_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ _05471_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _07168_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__xnor2_1
X_18901_ rbzero.pov.spi_buffer\[58\] rbzero.pov.ready_buffer\[58\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11236_ rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__inv_2
XFILLER_136_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19881_ net55 rbzero.pov.sclk_buffer\[0\] _09734_ vssd1 vssd1 vccd1 vccd1 _03553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18832_ rbzero.pov.spi_buffer\[25\] rbzero.pov.ready_buffer\[25\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02996_ sky130_fd_sc_hd__mux2_1
X_11167_ _04385_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18763_ _02952_ _02956_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__nor2_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _08528_ _08571_ _09069_ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__a21oi_1
X_11098_ rbzero.tex_b0\[54\] rbzero.tex_b0\[53\] _04340_ vssd1 vssd1 vccd1 vccd1 _04349_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17714_ _09519_ _09890_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__and2_1
XFILLER_76_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14926_ _08036_ _08063_ _08064_ _08061_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__o211a_1
X_18694_ _02887_ _02888_ _02892_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__or3_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17645_ _01927_ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__xnor2_1
X_14857_ rbzero.wall_tracer.stepDistY\[4\] _08012_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08013_ sky130_fd_sc_hd__mux2_1
XFILLER_1_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _06937_ _06938_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__xnor2_1
X_17576_ _01864_ _01866_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__o21ai_4
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14788_ _06581_ _07952_ _07866_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__o21a_1
XFILLER_189_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20303__168 clknet_1_0__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__inv_2
XFILLER_189_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19315_ rbzero.spi_registers.got_new_leak _03095_ vssd1 vssd1 vccd1 vccd1 _03272_
+ sky130_fd_sc_hd__and2_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16527_ _09498_ _09615_ _09616_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13739_ _06906_ _06905_ _06909_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__o21bai_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19246_ rbzero.spi_registers.new_texadd\[2\]\[18\] _03221_ _03232_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__o211a_1
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ _09547_ _09548_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15409_ _08500_ _08501_ _08503_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__a21bo_1
X_16389_ _09457_ _09459_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__or2_1
XFILLER_118_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19177_ rbzero.spi_registers.texadd1\[13\] _03189_ vssd1 vssd1 vccd1 vccd1 _03193_
+ sky130_fd_sc_hd__or2_1
XFILLER_145_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18128_ _02400_ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__o21a_1
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18059_ _02334_ _02342_ _02343_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__and3_1
XFILLER_28_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21070_ clknet_leaf_81_i_clk _00659_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ rbzero.pov.ready_buffer\[33\] _03656_ _03659_ _03630_ vssd1 vssd1 vccd1 vccd1
+ _01197_ sky130_fd_sc_hd__o211a_1
XFILLER_99_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21972_ net498 _01561_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ clknet_leaf_55_i_clk _00512_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20854_ clknet_leaf_51_i_clk _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20785_ gpout3.clk_div\[0\] net63 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__nor2_1
XFILLER_161_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21406_ clknet_leaf_28_i_clk _00995_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21337_ clknet_leaf_22_i_clk _00926_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ rbzero.tex_r1\[49\] _04981_ _05236_ _04918_ vssd1 vssd1 vccd1 vccd1 _05259_
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21268_ clknet_leaf_27_i_clk _00857_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11021_ rbzero.tex_b1\[26\] rbzero.tex_b1\[27\] _04303_ vssd1 vssd1 vccd1 vccd1 _04309_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21199_ clknet_leaf_29_i_clk _00788_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _08841_ _08842_ _08854_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__a21o_1
XFILLER_79_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ rbzero.map_overlay.i_mapdx\[1\] _06117_ _06120_ rbzero.map_overlay.i_mapdx\[2\]
+ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__o221a_1
XFILLER_79_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03806_ clknet_0__03806_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03806_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _05089_ _05097_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__nor2_4
X_14711_ _06580_ _07876_ _07877_ _07880_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__o31a_1
XFILLER_206_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _08770_ _08769_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__xor2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _09542_ _09560_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nor2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14642_ _06580_ _07807_ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__o21ai_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _05019_ _05041_ _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a21o_1
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _04195_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17361_ _10261_ _10264_ _10377_ _10378_ vssd1 vssd1 vccd1 vccd1 _10379_ sky130_fd_sc_hd__o211a_1
X_14573_ _07711_ _07716_ _07742_ _07743_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__and4_1
XFILLER_198_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11785_ _04947_ _04972_ _04974_ _04919_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__o211a_1
XFILLER_198_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19100_ rbzero.spi_registers.texadd0\[4\] _03143_ vssd1 vssd1 vccd1 vccd1 _03149_
+ sky130_fd_sc_hd__or2_1
XFILLER_207_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16312_ _09386_ _09403_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13524_ _06625_ _06635_ _06589_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17292_ _10203_ _10212_ _10310_ vssd1 vssd1 vccd1 vccd1 _10311_ sky130_fd_sc_hd__a21oi_1
X_10736_ _04159_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16243_ _09333_ _09334_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__and2_1
X_19031_ rbzero.map_overlay.i_otherx\[4\] _03101_ vssd1 vssd1 vccd1 vccd1 _03107_
+ sky130_fd_sc_hd__or2_1
XFILLER_186_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13455_ _06624_ _06625_ _06589_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _04121_ vssd1 vssd1 vccd1 vccd1 _04123_
+ sky130_fd_sc_hd__mux2_1
X_12406_ _04902_ _05586_ _05590_ _04823_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__o31a_1
XFILLER_185_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16174_ _09265_ _09266_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__xor2_1
XFILLER_177_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13386_ _06413_ _06487_ _06533_ _06465_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a221o_1
X_10598_ _04086_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15125_ rbzero.debug_overlay.playerY\[-6\] vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__inv_2
XFILLER_86_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12337_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _04907_ vssd1 vssd1 vccd1 vccd1 _05523_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15056_ _08150_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__clkbuf_4
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19933_ rbzero.debug_overlay.playerX\[1\] _03587_ _03582_ vssd1 vssd1 vccd1 vccd1
+ _03592_ sky130_fd_sc_hd__a21o_1
X_12268_ _04902_ _05441_ _05445_ _04823_ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a311o_1
XFILLER_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14007_ _06540_ _06942_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__or3_1
X_11219_ _04413_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__nor2_2
XFILLER_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19864_ _03544_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
X_12199_ rbzero.tex_g1\[13\] _04905_ _05186_ _04940_ vssd1 vssd1 vccd1 vccd1 _05386_
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03464_ _03464_ vssd1 vssd1 vccd1 vccd1 clknet_0__03464_ sky130_fd_sc_hd__clkbuf_16
X_18815_ rbzero.pov.spi_buffer\[17\] rbzero.pov.ready_buffer\[17\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
X_20383__240 clknet_1_1__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__inv_2
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19795_ _03508_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ _02935_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nor3_1
XFILLER_97_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _09051_ _09052_ _08357_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__a21o_2
XFILLER_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ _08036_ _08051_ _08052_ _01633_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__o211a_1
X_18677_ _02876_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__xnor2_1
X_15889_ _08898_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__inv_2
XFILLER_52_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17628_ _01813_ _01825_ _01823_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a21o_1
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17559_ _01848_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__xor2_1
XFILLER_177_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19229_ rbzero.spi_registers.new_texadd\[2\]\[10\] _03221_ _03223_ _03213_ vssd1
+ vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__o211a_1
XFILLER_164_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19669__49 clknet_1_0__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21122_ clknet_leaf_90_i_clk _00711_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20466__315 clknet_1_0__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__inv_2
XFILLER_120_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21053_ clknet_leaf_12_i_clk _00642_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20004_ rbzero.pov.ready_buffer\[56\] _03586_ _03644_ _03645_ _03617_ vssd1 vssd1
+ vccd1 vccd1 _03646_ sky130_fd_sc_hd__o221a_1
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ net481 _01544_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ clknet_leaf_36_i_clk _00495_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_203_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ net412 _01475_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ clknet_leaf_66_i_clk _00426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ _04756_ _04757_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__nand3_1
X_20768_ rbzero.wall_tracer.rayAddendY\[-8\] _02606_ _02557_ _03952_ vssd1 vssd1 vccd1
+ vccd1 _01652_ sky130_fd_sc_hd__a22o_1
XFILLER_35_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ rbzero.tex_r1\[5\] rbzero.tex_r1\[6\] _04035_ vssd1 vssd1 vccd1 vccd1 _04044_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20699_ rbzero.traced_texa\[8\] rbzero.texV\[8\] _03910_ vssd1 vssd1 vccd1 vccd1
+ _03915_ sky130_fd_sc_hd__a21o_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13240_ _06324_ _06328_ _06410_ _06322_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__a31oi_4
X_10452_ rbzero.tex_r1\[38\] rbzero.tex_r1\[39\] _04002_ vssd1 vssd1 vccd1 vccd1 _04008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ rbzero.wall_tracer.visualWallDist\[1\] _04427_ vssd1 vssd1 vccd1 vccd1 _06342_
+ sky130_fd_sc_hd__or2_1
XFILLER_108_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12122_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _04932_ vssd1 vssd1 vccd1 vccd1 _05310_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20332__194 clknet_1_0__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__inv_2
XFILLER_151_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16930_ _09940_ _09951_ vssd1 vssd1 vccd1 vccd1 _09952_ sky130_fd_sc_hd__xnor2_1
X_12053_ rbzero.tex_r1\[32\] _04982_ _04910_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_
+ sky130_fd_sc_hd__a31o_1
XFILLER_85_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ rbzero.tex_b1\[34\] rbzero.tex_b1\[35\] _04292_ vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16861_ _09874_ _09876_ _09875_ vssd1 vssd1 vccd1 vccd1 _09884_ sky130_fd_sc_hd__a21boi_1
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18600_ _02798_ _02799_ _02806_ _04434_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15812_ _08899_ _08895_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__nand2_1
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19580_ _03418_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__clkbuf_1
X_16792_ _09822_ _09108_ vssd1 vssd1 vccd1 vccd1 _09823_ sky130_fd_sc_hd__nand2_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18531_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__nor2_1
X_15743_ _08516_ _08344_ _08827_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__nor3_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ rbzero.debug_overlay.playerX\[4\] _06129_ _06130_ rbzero.debug_overlay.playerY\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__o22ai_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11906_ _05093_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18462_ _02598_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _02688_
+ sky130_fd_sc_hd__or2_1
XFILLER_179_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15674_ _08767_ _08768_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__xor2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _06060_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _10318_ _01705_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__xnor2_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ rbzero.row_render.side vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__inv_2
XFILLER_18_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14625_ _07626_ _07673_ _07793_ _07795_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__a22o_1
X_18393_ _02598_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02624_
+ sky130_fd_sc_hd__nand2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _10361_ _10362_ vssd1 vssd1 vccd1 vccd1 _10363_ sky130_fd_sc_hd__nand2_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14556_ _06959_ _07209_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__nor2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _04823_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__buf_6
XFILLER_147_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10719_ _04150_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13507_ _06469_ _06568_ _06594_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and3_1
X_17275_ _08666_ _09131_ vssd1 vssd1 vccd1 vccd1 _10294_ sky130_fd_sc_hd__nor2_1
X_14487_ _07654_ _07656_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11699_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__buf_6
XFILLER_186_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19014_ _05270_ _03091_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__and3_1
X_16226_ _09305_ _09318_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__xnor2_2
X_13438_ _06607_ _06608_ _06576_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__mux2_1
XFILLER_127_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20415__269 clknet_1_1__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__inv_2
X_16157_ _09248_ _09249_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _06379_ _06515_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__nor2_8
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04634_ _04634_ vssd1 vssd1 vccd1 vccd1 clknet_0__04634_ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15108_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__o21ai_1
X_16088_ _09177_ _09180_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__nor2_1
X_15039_ _08135_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__buf_6
X_19916_ _03212_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ rbzero.pov.spi_buffer\[60\] rbzero.pov.spi_buffer\[61\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03536_ sky130_fd_sc_hd__mux2_1
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19778_ _03499_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
X_20309__174 clknet_1_1__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__inv_2
XFILLER_209_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18729_ _04434_ _02924_ _02925_ _02889_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a22o_1
XFILLER_97_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21740_ net266 _01329_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21671_ clknet_leaf_25_i_clk _01260_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20622_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03850_
+ sky130_fd_sc_hd__nand2_1
XFILLER_189_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ clknet_leaf_70_i_clk _00694_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21036_ clknet_leaf_80_i_clk _00625_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12740_ net32 net33 vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__and2b_1
X_21938_ net464 _01527_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
X_20520__364 clknet_1_0__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__inv_2
XFILLER_167_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12671_ net51 _05842_ _05843_ net40 _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a221o_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21869_ net395 _01458_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _07045_ _07204_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__nor2_1
X_11622_ _04792_ _04806_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__nor3_4
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15390_ _08445_ _08484_ _08459_ _08474_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__a31oi_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14341_ _07503_ _07511_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11553_ _04698_ _04647_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ _03979_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__clkbuf_4
X_17060_ _10079_ _10080_ _09967_ _09965_ vssd1 vssd1 vccd1 vccd1 _10081_ sky130_fd_sc_hd__a22oi_2
XFILLER_183_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14272_ _07159_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__nor2_1
XFILLER_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ rbzero.debug_overlay.playerX\[2\] vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__clkinv_2
XFILLER_171_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16011_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerX\[-7\] _08138_
+ vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _06310_ _06312_ _06316_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__o21ai_1
X_10435_ rbzero.tex_r1\[46\] rbzero.tex_r1\[47\] _03991_ vssd1 vssd1 vccd1 vccd1 _03999_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _05996_ _05998_ _06029_ _06031_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a31o_1
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _05047_ _05266_ _05268_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__o31a_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _02248_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__and2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13085_ rbzero.trace_state\[0\] _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__or2_2
X_16913_ _09933_ _09934_ vssd1 vssd1 vccd1 vccd1 _09935_ sky130_fd_sc_hd__nor2_1
X_12036_ _04955_ _05211_ _05215_ _04887_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a311o_1
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17893_ _02179_ _02180_ _06105_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a21oi_1
X_19632_ rbzero.pov.spi_counter\[3\] _03448_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__nand2_1
X_16844_ _06104_ _09868_ vssd1 vssd1 vccd1 vccd1 _09869_ sky130_fd_sc_hd__nand2_1
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19563_ rbzero.spi_registers.new_texadd\[0\]\[23\] rbzero.spi_registers.spi_buffer\[23\]
+ _03380_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XFILLER_207_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775_ _06189_ _09786_ _09807_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a21oi_1
X_13987_ _07157_ _07053_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__xnor2_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _04674_ _02729_ _08124_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
X_15726_ _08766_ _08817_ _08820_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__o21a_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ rbzero.spi_registers.new_mapd\[11\] rbzero.spi_registers.spi_buffer\[11\]
+ _03361_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__mux2_1
X_12938_ rbzero.debug_overlay.playerY\[5\] vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__inv_2
XFILLER_179_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20495__341 clknet_1_1__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__inv_2
X_18445_ _02653_ _02670_ _02671_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__or3_1
XFILLER_181_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15657_ _08748_ _08750_ _08751_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__a21o_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _06042_ _06043_ _06025_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__or3b_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14608_ _07763_ _07766_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__nor2_1
X_18376_ _02596_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02608_
+ sky130_fd_sc_hd__and2_1
X_15588_ _08287_ _08336_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__nor2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327_ _10096_ _10219_ _10221_ vssd1 vssd1 vccd1 vccd1 _10346_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14539_ _07645_ _07665_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ _09525_ _09362_ _10276_ vssd1 vssd1 vccd1 vccd1 _10277_ sky130_fd_sc_hd__o21a_1
XFILLER_31_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16209_ _08434_ _09037_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__nor2_1
X_17189_ _10207_ _10208_ vssd1 vssd1 vccd1 vccd1 _10209_ sky130_fd_sc_hd__nand2_1
XFILLER_127_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21723_ net249 _01312_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21654_ clknet_leaf_43_i_clk _01243_ vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_200_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20605_ _03830_ _03832_ _03831_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21bai_1
XFILLER_177_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21585_ clknet_leaf_91_i_clk _01174_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_77 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_77/HI o_rgb[2] sky130_fd_sc_hd__conb_1
XFILLER_71_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_88 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_88/HI o_rgb[17] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_99 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_99/HI zeros[6] sky130_fd_sc_hd__conb_1
XFILLER_165_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22068_ clknet_leaf_40_i_clk _01657_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13910_ _07076_ _07077_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__a21oi_1
X_21019_ clknet_leaf_74_i_clk _00608_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14890_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1 vccd1 vccd1 _08039_
+ sky130_fd_sc_hd__inv_2
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13841_ _06973_ _07009_ _07010_ _06971_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__a22o_1
X_20444__295 clknet_1_1__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__inv_2
XFILLER_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _09522_ _09649_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__xor2_1
X_13772_ _06682_ _06693_ _06941_ _06942_ _06754_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__o32a_1
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10984_ _04289_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15511_ _08597_ _08593_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__or2b_1
X_12723_ _05889_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__inv_2
X_16491_ _09580_ _09581_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__and2b_1
XFILLER_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18230_ rbzero.spi_registers.spi_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__clkbuf_4
X_15442_ _08150_ _08335_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__nor2_1
X_12654_ net23 vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__inv_2
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _04760_ _04793_ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a21o_1
XFILLER_129_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18161_ _02429_ _02430_ _02424_ _02427_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a211oi_1
XFILLER_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15373_ _08459_ _08467_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__xnor2_1
X_12585_ net19 vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__inv_2
XFILLER_157_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _09866_ _10131_ _10132_ vssd1 vssd1 vccd1 vccd1 _10133_ sky130_fd_sc_hd__or3b_1
X_14324_ _07486_ _07487_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__nand2_1
X_11536_ rbzero.map_overlay.i_mapdx\[5\] _04725_ _04720_ vssd1 vssd1 vccd1 vccd1 _04726_
+ sky130_fd_sc_hd__o21a_1
X_18092_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__nor2_1
XFILLER_102_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03781_ _03781_ vssd1 vssd1 vccd1 vccd1 clknet_0__03781_ sky130_fd_sc_hd__clkbuf_16
X_17043_ _10062_ _10063_ vssd1 vssd1 vccd1 vccd1 _10064_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ _07303_ _06807_ _06808_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__and3b_1
X_11467_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__clkbuf_4
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _06375_ _06376_ _06323_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__mux2_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10418_ rbzero.tex_r1\[54\] rbzero.tex_r1\[55\] _03980_ vssd1 vssd1 vccd1 vccd1 _03990_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186_ _07327_ _07356_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11398_ _04509_ _04481_ _04507_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__and3_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _06292_ _06294_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__and2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ rbzero.spi_registers.spi_cmd\[3\] _02475_ _03078_ vssd1 vssd1 vccd1 vccd1
+ _03082_ sky130_fd_sc_hd__mux2_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _02226_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__and2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ rbzero.map_overlay.i_othery\[2\] _06086_ _06107_ rbzero.map_overlay.i_othery\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__o22a_1
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ rbzero.tex_r1\[22\] _05182_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or2_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17876_ _01994_ _02069_ _02164_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a21oi_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19615_ _03100_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__nand2_1
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16827_ _06183_ _09786_ _09853_ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19546_ _03401_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16758_ _09790_ _09793_ vssd1 vssd1 vccd1 vccd1 _09794_ sky130_fd_sc_hd__xor2_1
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15709_ _08746_ _08784_ _08800_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__nand3_1
XFILLER_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19477_ _03365_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16689_ rbzero.row_render.texu\[1\] _09752_ _09754_ rbzero.texu_hot\[1\] vssd1 vssd1
+ vccd1 vccd1 _00495_ sky130_fd_sc_hd__a22o_1
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18428_ _02655_ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__nand2_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__inv_2
XFILLER_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21370_ clknet_leaf_12_i_clk _00959_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20183_ rbzero.spi_registers.new_texadd\[3\]\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__mux2_1
XFILLER_153_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21706_ net232 _01295_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21637_ clknet_leaf_82_i_clk _01226_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _05029_ _05554_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 _05555_
+ sky130_fd_sc_hd__or3b_1
XFILLER_201_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21568_ clknet_leaf_93_i_clk _01157_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11321_ _04477_ _04510_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21499_ clknet_leaf_98_i_clk _01088_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14040_ _07205_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__and2b_1
X_11252_ _04444_ _04441_ _04435_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a21bo_1
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11183_ _04393_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15991_ _08568_ _09074_ _09085_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__a21oi_4
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17730_ _01894_ _01907_ _01905_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a21oi_1
X_14942_ rbzero.wall_tracer.visualWallDist\[3\] _08046_ vssd1 vssd1 vccd1 vccd1 _08076_
+ sky130_fd_sc_hd__or2_1
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17661_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__nor2_1
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14873_ _06470_ _06598_ _07871_ _07989_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__a31o_1
XFILLER_36_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19400_ _03322_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
X_16612_ _09572_ _09573_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__nor2_1
X_13824_ _06757_ _06854_ _06985_ _06681_ _06693_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a32o_1
X_17592_ _01827_ _01805_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__or2b_1
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19331_ rbzero.color_sky\[0\] _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__a21o_1
X_16543_ _09625_ _09632_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__xnor2_1
X_10967_ _04280_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
X_13755_ _06919_ _06924_ _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__or3_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ net31 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__inv_2
X_19262_ rbzero.spi_registers.texadd3\[0\] _03242_ vssd1 vssd1 vccd1 vccd1 _03243_
+ sky130_fd_sc_hd__or2_1
XFILLER_203_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16474_ _08027_ _09563_ _08029_ vssd1 vssd1 vccd1 vccd1 _09565_ sky130_fd_sc_hd__o21ai_1
X_10898_ _04244_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
X_13686_ _06856_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__clkbuf_2
XFILLER_204_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18213_ _02475_ _02476_ _04052_ rbzero.spi_registers.spi_done vssd1 vssd1 vccd1 vccd1
+ _02477_ sky130_fd_sc_hd__or4b_4
X_15425_ _08517_ _08518_ _08519_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__a21bo_1
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ _05799_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nand2_1
X_19193_ rbzero.spi_registers.new_texadd\[1\]\[20\] _03173_ _03201_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__o211a_1
XFILLER_19_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03802_ clknet_0__03802_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03802_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18144_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__nand2_1
X_12568_ net11 _05704_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__nand2_1
XFILLER_106_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15356_ _08000_ _08425_ _08006_ vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19704__81 clknet_1_0__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14307_ _07445_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__and2_1
X_11519_ _04656_ rbzero.map_overlay.i_othery\[2\] vssd1 vssd1 vccd1 vccd1 _04709_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18075_ _02341_ _02356_ _02357_ _02337_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__o31a_1
XFILLER_117_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15287_ _08381_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12499_ _03975_ _04420_ _05646_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__mux2_1
XFILLER_116_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _10045_ _10046_ vssd1 vssd1 vccd1 vccd1 _10047_ sky130_fd_sc_hd__xor2_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14238_ _07395_ _07407_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and3_1
XFILLER_172_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14169_ _07336_ _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__nand2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ rbzero.spi_registers.spi_buffer\[19\] rbzero.spi_registers.spi_buffer\[18\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ rbzero.wall_tracer.visualWallDist\[8\] _01699_ vssd1 vssd1 vccd1 vccd1 _02216_
+ sky130_fd_sc_hd__nand2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17859_ _02146_ _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__nor2_1
XFILLER_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20870_ clknet_leaf_43_i_clk _00459_ vssd1 vssd1 vccd1 vccd1 reg_rgb\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19529_ _03392_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_i_clk clknet_1_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1_1_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21422_ clknet_leaf_4_i_clk _01011_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21353_ clknet_leaf_35_i_clk _00942_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vshift
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21284_ clknet_leaf_2_i_clk _00873_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20235_ clknet_1_0__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__buf_1
XFILLER_162_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20166_ _05653_ _03747_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nand2_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20097_ _03084_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__buf_4
XFILLER_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _05059_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ rbzero.tex_g0\[58\] rbzero.tex_g0\[57\] _04203_ vssd1 vssd1 vccd1 vccd1 _04204_
+ sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20999_ clknet_leaf_0_i_clk _00588_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ rbzero.tex_g1\[26\] rbzero.tex_g1\[27\] _04166_ vssd1 vssd1 vccd1 vccd1 _04168_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13540_ _06547_ _06579_ _06633_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__o21ai_1
XFILLER_186_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _06508_ _06482_ _06565_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__mux2_1
XFILLER_197_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ rbzero.tex_g1\[58\] rbzero.tex_g1\[59\] _04046_ vssd1 vssd1 vccd1 vccd1 _04131_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15210_ _08152_ _08304_ _08166_ _08171_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__o22ai_2
X_12422_ _04922_ _05604_ _05605_ _05606_ _04940_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__o221a_1
XFILLER_205_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _09280_ _09282_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__xor2_1
XFILLER_205_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15141_ _08228_ _08235_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__nor2_1
X_12353_ _04823_ _05514_ _05522_ _05538_ _04832_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a311o_1
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ rbzero.texu_hot\[0\] _04494_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nand3_1
X_15072_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] _04463_
+ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__mux2_1
X_12284_ reg_rgb\[15\] _05470_ _05058_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__mux2_2
XFILLER_114_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14023_ _07192_ _07193_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__nand2_1
XFILLER_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18900_ _03031_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
X_11235_ rbzero.trace_state\[1\] rbzero.trace_state\[0\] vssd1 vssd1 vccd1 vccd1 _04430_
+ sky130_fd_sc_hd__or2_2
X_19880_ _03552_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _02995_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
X_11166_ rbzero.tex_b0\[22\] rbzero.tex_b0\[21\] _04384_ vssd1 vssd1 vccd1 vccd1 _04385_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18762_ rbzero.spi_registers.spi_counter\[2\] _02955_ vssd1 vssd1 vccd1 vccd1 _02956_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15974_ _08495_ _08527_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__and2b_1
X_11097_ _04348_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17713_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__xor2_1
X_14925_ rbzero.wall_tracer.visualWallDist\[-2\] _08047_ vssd1 vssd1 vccd1 vccd1 _08064_
+ sky130_fd_sc_hd__or2_1
X_18693_ _02887_ _02888_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__o21ai_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _01933_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__nor2_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14856_ _08011_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__buf_2
XFILLER_1_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13807_ _06726_ _06785_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or3_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _01864_ _01866_ _01757_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14787_ _07950_ _07951_ _06574_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__mux2_1
X_11999_ rbzero.tex_r1\[12\] _04906_ _05181_ _05184_ _05187_ vssd1 vssd1 vccd1 vccd1
+ _05188_ sky130_fd_sc_hd__a311o_1
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19314_ rbzero.spi_registers.got_new_leak _03097_ vssd1 vssd1 vccd1 vccd1 _03271_
+ sky130_fd_sc_hd__nand2_2
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16526_ _09005_ _09252_ _09243_ _08952_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__o22a_1
XFILLER_182_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ _06901_ _06903_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19245_ rbzero.spi_registers.texadd2\[18\] _03222_ vssd1 vssd1 vccd1 vccd1 _03232_
+ sky130_fd_sc_hd__or2_1
X_16457_ _09044_ _09046_ _08369_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ _06834_ _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _08042_ _08428_ _08502_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__or3_1
X_19176_ rbzero.spi_registers.new_texadd\[1\]\[12\] _03188_ _03192_ _03184_ vssd1
+ vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__o211a_1
X_16388_ _09344_ _09346_ _09466_ _09478_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__a31oi_4
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18127_ _02400_ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__nor3_1
X_15339_ _08228_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18058_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__nand2_1
XFILLER_67_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17009_ _09146_ _09242_ _09363_ _09005_ vssd1 vssd1 vccd1 vccd1 _10030_ sky130_fd_sc_hd__o22a_1
XFILLER_160_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ rbzero.debug_overlay.facingX\[-9\] _03658_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__or2_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21971_ net497 _01560_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20922_ clknet_leaf_56_i_clk _00511_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ clknet_leaf_51_i_clk _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20784_ _03962_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20278__146 clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__inv_2
XFILLER_35_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21405_ clknet_leaf_32_i_clk _00994_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21336_ clknet_leaf_9_i_clk _00925_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21267_ clknet_leaf_27_i_clk _00856_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11020_ _04308_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21198_ clknet_leaf_28_i_clk _00787_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20149_ _05648_ _03093_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2_1
XFILLER_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03805_ clknet_0__03805_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03805_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ rbzero.map_overlay.i_mapdx\[3\] rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1
+ _06147_ sky130_fd_sc_hd__xnor2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14710_ _06580_ _07879_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__nand2_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11922_ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__buf_4
X_15690_ _08738_ _08740_ _08739_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__a21o_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14641_ _06580_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__nand2_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _05027_ _05042_ _05017_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a21o_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ rbzero.tex_g1\[1\] rbzero.tex_g1\[2\] _04188_ vssd1 vssd1 vccd1 vccd1 _04195_
+ sky130_fd_sc_hd__mux2_1
X_17360_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _10378_ sky130_fd_sc_hd__or2_1
XFILLER_14_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11784_ _04934_ _04973_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or2_1
X_14572_ _07710_ _07709_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__xor2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16311_ _09392_ _09402_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__xor2_1
XFILLER_201_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _06644_ _06653_ _06641_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__mux2_1
X_17291_ _10206_ _10211_ vssd1 vssd1 vccd1 vccd1 _10310_ sky130_fd_sc_hd__and2b_1
X_10735_ rbzero.tex_g1\[34\] rbzero.tex_g1\[35\] _04155_ vssd1 vssd1 vccd1 vccd1 _04159_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ rbzero.spi_registers.new_other\[9\] _03098_ _03106_ _03103_ vssd1 vssd1 vccd1
+ vccd1 _00759_ sky130_fd_sc_hd__o211a_1
X_16242_ _09333_ _09334_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__nor2_1
X_10666_ _04122_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13454_ _06458_ _06465_ _06578_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__mux2_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ _04922_ _05587_ _05589_ _04940_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__o211a_1
X_16173_ _09081_ _09136_ _09075_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__or3b_1
X_13385_ _06430_ _06432_ _06555_ _06547_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__a22o_1
X_10597_ rbzero.tex_r0\[36\] rbzero.tex_r0\[35\] _04077_ vssd1 vssd1 vccd1 vccd1 _04086_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ _08217_ rbzero.debug_overlay.playerX\[-6\] _08218_ vssd1 vssd1 vccd1 vccd1
+ _08219_ sky130_fd_sc_hd__mux2_1
X_12336_ _04953_ _05517_ _05521_ _04812_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a211o_1
XFILLER_115_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15055_ rbzero.wall_tracer.visualWallDist\[1\] _08149_ vssd1 vssd1 vccd1 vccd1 _08150_
+ sky130_fd_sc_hd__nand2_2
X_12267_ _05447_ _05449_ _05451_ _05453_ _04889_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__o221a_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19932_ rbzero.debug_overlay.playerX\[1\] _03587_ vssd1 vssd1 vccd1 vccd1 _03591_
+ sky130_fd_sc_hd__nor2_1
X_14006_ _06710_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__xnor2_1
X_11218_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__inv_4
X_19863_ rbzero.pov.spi_buffer\[68\] rbzero.pov.spi_buffer\[69\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03544_ sky130_fd_sc_hd__mux2_1
X_12198_ rbzero.tex_g1\[15\] _04910_ _05384_ _04912_ vssd1 vssd1 vccd1 vccd1 _05385_
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03463_ _03463_ vssd1 vssd1 vccd1 vccd1 clknet_0__03463_ sky130_fd_sc_hd__clkbuf_16
X_11149_ rbzero.tex_b0\[30\] rbzero.tex_b0\[29\] _04373_ vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__mux2_1
X_18814_ _02986_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19794_ rbzero.pov.spi_buffer\[35\] rbzero.pov.spi_buffer\[36\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18745_ _02939_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__nand2_1
XFILLER_49_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15957_ rbzero.wall_tracer.stepDistY\[5\] _08338_ vssd1 vssd1 vccd1 vccd1 _09052_
+ sky130_fd_sc_hd__nand2_1
XFILLER_23_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14908_ rbzero.wall_tracer.visualWallDist\[-7\] _08047_ vssd1 vssd1 vccd1 vccd1 _08052_
+ sky130_fd_sc_hd__or2_1
XFILLER_209_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18676_ _02860_ _02866_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nand2_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _08971_ _08982_ _08978_ _08979_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17627_ _01881_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14839_ _07997_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17558_ _01715_ _01737_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16509_ rbzero.texu_hot\[4\] _08145_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__or2_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17489_ _09519_ _09363_ _10276_ _01666_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__o31a_1
XFILLER_34_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19228_ rbzero.spi_registers.texadd2\[10\] _03222_ vssd1 vssd1 vccd1 vccd1 _03223_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19159_ rbzero.spi_registers.new_texadd\[1\]\[5\] _03174_ _03182_ _03169_ vssd1 vssd1
+ vccd1 vccd1 _00812_ sky130_fd_sc_hd__o211a_1
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21121_ clknet_leaf_91_i_clk _00710_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21052_ clknet_leaf_12_i_clk _00641_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20003_ rbzero.debug_overlay.playerY\[3\] _03640_ _03116_ vssd1 vssd1 vccd1 vccd1
+ _03645_ sky130_fd_sc_hd__a21o_1
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ net480 _01543_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20905_ clknet_leaf_20_i_clk _00494_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_199_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21885_ net411 _01474_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20836_ clknet_leaf_60_i_clk _00425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20767_ _02747_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ _04043_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20698_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03914_
+ sky130_fd_sc_hd__nand2_1
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ _04007_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13170_ _06339_ _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20548__9 clknet_1_1__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12121_ _04923_ _05306_ _05307_ _05308_ _04941_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__o221a_1
X_21319_ clknet_leaf_31_i_clk _00908_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ rbzero.tex_r1\[33\] _04981_ _05236_ _04918_ vssd1 vssd1 vccd1 vccd1 _05241_
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11003_ _04299_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16860_ _09881_ _09882_ vssd1 vssd1 vccd1 vccd1 _09883_ sky130_fd_sc_hd__or2_1
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ _08867_ _08902_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__xnor2_1
X_16791_ _06103_ vssd1 vssd1 vccd1 vccd1 _09822_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18530_ _02742_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__clkbuf_1
X_15742_ _08799_ _08836_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__nand2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__clkinv_2
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ rbzero.wall_tracer.rayAddendX\[8\] _02527_ _02680_ _02687_ vssd1 vssd1 vccd1
+ vccd1 _00609_ sky130_fd_sc_hd__o22a_1
X_11905_ _05075_ _05081_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nand2_1
X_15673_ _08213_ _08269_ _08274_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__or3_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12885_ _06013_ _06016_ _06011_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a21o_1
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _08814_ _09677_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__nor2_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _07626_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__xnor2_1
X_11836_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__inv_2
X_18392_ _02557_ _02612_ _02613_ _02623_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a31o_1
XFILLER_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _10271_ _10360_ vssd1 vssd1 vccd1 vccd1 _10362_ sky130_fd_sc_hd__or2_1
XFILLER_198_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14555_ _07693_ _07697_ _07695_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__o21ai_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _04903_ _04921_ _04938_ _04956_ _04887_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__o311a_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__05820_ _05820_ vssd1 vssd1 vccd1 vccd1 clknet_0__05820_ sky130_fd_sc_hd__clkbuf_16
X_13506_ _06641_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__or2_1
XFILLER_187_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17274_ _10291_ _10292_ vssd1 vssd1 vccd1 vccd1 _10293_ sky130_fd_sc_hd__nand2_1
X_10718_ rbzero.tex_g1\[42\] rbzero.tex_g1\[43\] _04144_ vssd1 vssd1 vccd1 vccd1 _04150_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14486_ _06729_ _07310_ _07655_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__nand3_1
XFILLER_105_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ _04792_ _04806_ _04811_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__or3_1
XFILLER_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19013_ _05644_ _09747_ _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__and3_1
X_16225_ _09313_ _09317_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__xor2_2
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13437_ _06451_ _06458_ _06565_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__mux2_1
X_10649_ _04113_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ _08296_ _08617_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__nor2_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13368_ _06494_ _06538_ _06535_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or3_4
XFILLER_177_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15107_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__or3_1
XFILLER_154_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12319_ _04812_ _05492_ _05496_ _05504_ _04886_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__o311a_1
X_16087_ _09177_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__and2_1
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13299_ _06469_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__clkbuf_4
X_15038_ _08134_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__buf_4
X_19915_ rbzero.pov.ready_buffer\[65\] _03438_ _03558_ _03577_ vssd1 vssd1 vccd1 vccd1
+ _03578_ sky130_fd_sc_hd__a211o_1
XFILLER_190_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _03535_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16989_ _09872_ _10010_ vssd1 vssd1 vccd1 vccd1 _10011_ sky130_fd_sc_hd__nand2_1
X_19777_ rbzero.pov.spi_buffer\[27\] rbzero.pov.spi_buffer\[28\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XFILLER_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18728_ _02794_ _02911_ _08134_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__o21a_1
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18659_ _05127_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02861_
+ sky130_fd_sc_hd__or2_1
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21670_ clknet_leaf_31_i_clk _01259_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20621_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03849_
+ sky130_fd_sc_hd__nor2_1
XFILLER_196_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20472__320 clknet_1_0__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__inv_2
XFILLER_178_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_191_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21104_ clknet_leaf_70_i_clk _00693_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21035_ clknet_leaf_80_i_clk _00624_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21937_ net463 _01526_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ net41 _05845_ _05847_ _05263_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a22o_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21868_ net394 _01457_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _04767_ _04791_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and2_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ clknet_leaf_63_i_clk _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21799_ net325 _01388_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ _07505_ _07510_ _07509_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__a21o_1
X_11552_ _04722_ _04729_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o21a_1
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10503_ _04034_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14271_ _07156_ _07158_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__and2_1
XFILLER_52_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__inv_2
XFILLER_11_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _08997_ _08999_ vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__xor2_4
XFILLER_155_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10434_ _03998_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13222_ _06350_ _06352_ _06356_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a211oi_4
XFILLER_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13153_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__buf_4
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _05278_ _05291_ _05292_ _04744_ _04703_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a221o_1
XFILLER_152_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17961_ _02152_ _02246_ _02247_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__nand3_1
XFILLER_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13084_ rbzero.trace_state\[1\] _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nand2_4
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16912_ _08166_ _08382_ vssd1 vssd1 vccd1 vccd1 _09934_ sky130_fd_sc_hd__nor2_1
X_12035_ _05217_ _05219_ _05221_ _05223_ _04903_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__o221a_1
X_17892_ _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__05938_ clknet_0__05938_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05938_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16843_ _09355_ _09466_ vssd1 vssd1 vccd1 vccd1 _09868_ sky130_fd_sc_hd__xnor2_4
X_19631_ _03448_ _03449_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__nor2_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ _03409_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__clkbuf_1
X_16774_ _09782_ _09804_ _09806_ vssd1 vssd1 vccd1 vccd1 _09807_ sky130_fd_sc_hd__and3_1
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13986_ _07054_ _07043_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__and2b_1
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18513_ _09768_ _09771_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__xnor2_1
X_15725_ _08818_ _08819_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__or2b_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19493_ _03373_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12937_ rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__clkbuf_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18444_ _02670_ _02671_ _02653_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__o21ai_1
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15656_ _08728_ _08747_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__nor2_1
XFILLER_2_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12868_ _06042_ _06043_ _06025_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__o21bai_2
XFILLER_178_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _07776_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11819_ _04907_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__buf_4
X_18375_ rbzero.wall_tracer.rayAddendX\[2\] _02527_ _02601_ _02607_ vssd1 vssd1 vccd1
+ vccd1 _00603_ sky130_fd_sc_hd__o22a_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15587_ _08265_ _08298_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__nor2_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _05958_ _05057_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__or2_1
XFILLER_18_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ _10096_ _10344_ vssd1 vssd1 vccd1 vccd1 _10345_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ _07682_ _07707_ _07708_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__a21oi_2
XFILLER_202_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _09520_ _09242_ vssd1 vssd1 vccd1 vccd1 _10276_ sky130_fd_sc_hd__or2_1
XFILLER_30_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14469_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__clkbuf_2
XFILLER_128_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16208_ _09289_ _09300_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__xor2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17188_ _08816_ _09677_ _09560_ _08889_ vssd1 vssd1 vccd1 vccd1 _10208_ sky130_fd_sc_hd__o22ai_1
XFILLER_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _09229_ _09231_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__nand2_1
XFILLER_89_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19829_ _03526_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20504__349 clknet_1_0__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__inv_2
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21722_ net248 _01311_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21653_ clknet_leaf_46_i_clk _01242_ vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20604_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03835_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_138_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21584_ clknet_leaf_91_i_clk _01173_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_78 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_78/HI o_rgb[3] sky130_fd_sc_hd__conb_1
XFILLER_181_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_89 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_89/HI o_rgb[18] sky130_fd_sc_hd__conb_1
XFILLER_193_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22067_ clknet_leaf_36_i_clk _01656_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21018_ clknet_leaf_74_i_clk _00607_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _06971_ _06973_ _07009_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__nand4_1
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ _06750_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__clkbuf_4
X_10983_ rbzero.tex_b1\[44\] rbzero.tex_b1\[45\] _04281_ vssd1 vssd1 vccd1 vccd1 _04289_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15510_ _08596_ _08594_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__or2b_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _04687_ _04653_ _05645_ _04642_ _05881_ _05889_ vssd1 vssd1 vccd1 vccd1 _05900_
+ sky130_fd_sc_hd__mux4_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16490_ _09578_ _09579_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__nand2_1
XFILLER_203_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ _08331_ _08337_ _08535_ _08326_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__o31a_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12653_ net26 _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18160_ _02424_ _02427_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__o211a_1
X_11604_ _04757_ _04759_ _04756_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15372_ _08461_ _08466_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__or2_1
X_12584_ _05763_ _05057_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__or2_1
XFILLER_129_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17111_ _10128_ _10129_ _10130_ vssd1 vssd1 vccd1 vccd1 _10132_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14323_ _07432_ _07489_ _07490_ _07493_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__o22a_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11535_ rbzero.map_overlay.i_mapdx\[3\] rbzero.map_overlay.i_mapdx\[2\] rbzero.map_overlay.i_mapdx\[1\]
+ rbzero.map_overlay.i_mapdx\[0\] vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__or4_1
X_18091_ _09845_ _02371_ _02340_ rbzero.wall_tracer.trackDistY\[-6\] vssd1 vssd1 vccd1
+ vccd1 _00555_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _09647_ _08620_ vssd1 vssd1 vccd1 vccd1 _10063_ sky130_fd_sc_hd__nor2_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03780_ _03780_ vssd1 vssd1 vccd1 vccd1 clknet_0__03780_ sky130_fd_sc_hd__clkbuf_16
X_14254_ _07423_ _07398_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__o21ai_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__clkbuf_4
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ rbzero.wall_tracer.visualWallDist\[-9\] _06066_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__mux2_1
X_10417_ _03989_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14185_ _07341_ _07355_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__xor2_1
X_11397_ _04578_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__clkbuf_4
XFILLER_178_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _06293_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nor2_1
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _03081_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _02227_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__xor2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _04708_ _06113_ _06121_ rbzero.map_overlay.i_othery\[4\] _06242_ vssd1 vssd1
+ vccd1 vccd1 _06243_ sky130_fd_sc_hd__a221o_1
XFILLER_39_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _04903_ _05188_ _05194_ _04958_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a311o_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17875_ _02066_ _02068_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__nor2_1
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19614_ net41 net40 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__or2_2
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16826_ _06105_ _09851_ _09852_ _09812_ vssd1 vssd1 vccd1 vccd1 _09853_ sky130_fd_sc_hd__o211a_1
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19545_ rbzero.spi_registers.new_texadd\[0\]\[14\] rbzero.spi_registers.spi_buffer\[14\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16757_ _09763_ _09791_ _09792_ vssd1 vssd1 vccd1 vccd1 _09793_ sky130_fd_sc_hd__or3_1
X_13969_ _07081_ _07131_ _07138_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nor3_1
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15708_ _08782_ _08802_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__nor2_1
XFILLER_146_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19476_ rbzero.spi_registers.new_mapd\[2\] _02483_ _03362_ vssd1 vssd1 vccd1 vccd1
+ _03365_ sky130_fd_sc_hd__mux2_1
X_16688_ rbzero.row_render.texu\[0\] _09752_ _09754_ rbzero.texu_hot\[0\] vssd1 vssd1
+ vccd1 vccd1 _00494_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15639_ _08200_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__clkbuf_4
X_18427_ _05106_ _02642_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__nand2_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _02577_ _02587_ _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__o21a_1
XFILLER_175_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ _10309_ _10327_ vssd1 vssd1 vccd1 vccd1 _10328_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18289_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__nor2_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20182_ _03757_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21705_ net231 _01294_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21636_ clknet_leaf_80_i_clk _01225_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_166_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21567_ clknet_leaf_93_i_clk _01156_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ _04473_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or2_1
XFILLER_10_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21498_ clknet_leaf_98_i_clk _01087_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__buf_2
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11182_ rbzero.tex_b0\[14\] rbzero.tex_b0\[13\] _04384_ vssd1 vssd1 vccd1 vccd1 _04393_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15990_ _09083_ _09084_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__nand2_1
XFILLER_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14941_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.trackDistX\[3\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__mux2_1
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17660_ _01838_ _01842_ _01839_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a21boi_1
X_14872_ _08024_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
X_16611_ _09676_ _09700_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13823_ _06790_ _06727_ _06993_ _06772_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__o22a_1
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17591_ _01826_ _01808_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__or2b_1
X_16542_ _09626_ _09631_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__xor2_1
X_19330_ rbzero.spi_registers.new_sky\[0\] rbzero.spi_registers.got_new_sky _03097_
+ _04409_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a31o_1
X_13754_ _06849_ _06923_ _06922_ _06914_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a211oi_1
X_10966_ rbzero.tex_b1\[52\] rbzero.tex_b1\[53\] _04270_ vssd1 vssd1 vccd1 vccd1 _04280_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12705_ _05881_ _05297_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nand2_1
X_19261_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__clkbuf_4
XFILLER_206_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16473_ _08027_ _08029_ _09563_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__or3_1
X_13685_ _06742_ _06743_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__and2_1
XFILLER_204_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10897_ rbzero.tex_g0\[22\] rbzero.tex_g0\[21\] _04237_ vssd1 vssd1 vccd1 vccd1 _04244_
+ sky130_fd_sc_hd__mux2_1
X_18212_ rbzero.spi_registers.spi_cmd\[3\] vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__inv_2
X_15424_ _08235_ _08246_ _08371_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__or3_1
XFILLER_203_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _05765_ _05770_ _05814_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__a31o_1
X_19192_ rbzero.spi_registers.texadd1\[20\] _03175_ vssd1 vssd1 vccd1 vccd1 _03201_
+ sky130_fd_sc_hd__or2_1
XFILLER_54_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03801_ clknet_0__03801_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03801_
+ sky130_fd_sc_hd__clkbuf_16
X_18143_ _10127_ _02416_ _02364_ rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1
+ vccd1 _00562_ sky130_fd_sc_hd__o2bb2a_1
X_15355_ _08449_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__buf_2
XFILLER_156_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12567_ _04454_ _05719_ net14 _05703_ _05717_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a2111oi_1
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14306_ _06720_ _07476_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__nor2_1
XFILLER_89_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18074_ _02353_ _02354_ _02355_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a21oi_1
X_11518_ rbzero.map_overlay.i_otherx\[1\] vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__inv_2
X_15286_ rbzero.wall_tracer.stepDistY\[-2\] _08168_ _08380_ vssd1 vssd1 vccd1 vccd1
+ _08381_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _03969_ gpout0.hpos\[1\] _04452_ _04628_ _05646_ net5 vssd1 vssd1 vccd1 vccd1
+ _05680_ sky130_fd_sc_hd__mux4_1
X_17025_ _09525_ _09252_ vssd1 vssd1 vccd1 vccd1 _10046_ sky130_fd_sc_hd__nor2_1
XFILLER_176_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14237_ _07404_ _07406_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__nand2_1
X_11449_ gpout0.hpos\[5\] _04638_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04639_
+ sky130_fd_sc_hd__o21a_1
XFILLER_98_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14168_ _07249_ _07337_ _07338_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__a21o_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__or2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _03072_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__clkbuf_1
X_14099_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__inv_2
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17927_ _02099_ _02113_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a21bo_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17858_ _02006_ _02018_ _02016_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a21oi_1
X_20427__280 clknet_1_0__leaf__03795_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__inv_2
XFILLER_39_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _06105_ _09836_ _09837_ _09812_ vssd1 vssd1 vccd1 vccd1 _09838_ sky130_fd_sc_hd__o211a_1
X_17789_ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__inv_2
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19528_ rbzero.spi_registers.new_texadd\[0\]\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__mux2_1
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19459_ _03355_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21421_ clknet_leaf_4_i_clk _01010_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21352_ clknet_leaf_35_i_clk _00941_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21283_ clknet_leaf_100_i_clk _00872_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20165_ _05653_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__or2_1
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ _02756_ _03655_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__nand2_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10820_ _04054_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ clknet_leaf_0_i_clk _00587_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10751_ _04167_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13470_ _06610_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__clkbuf_4
X_10682_ _04130_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ rbzero.tex_b1\[2\] _04909_ _04981_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a21o_1
X_21619_ clknet_leaf_87_i_clk _01208_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
X_20255__125 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__inv_2
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15140_ _08234_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__clkbuf_4
X_12352_ _04812_ _05529_ _05537_ _04886_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__o211a_1
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ rbzero.spi_registers.texadd0\[6\] _04466_ vssd1 vssd1 vccd1 vccd1 _04495_
+ sky130_fd_sc_hd__or2_1
X_15071_ _08165_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12283_ rbzero.trace_state\[3\] _04635_ _05056_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_
+ sky130_fd_sc_hd__o211a_2
XFILLER_5_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14022_ _07181_ _07191_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nand2_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11234_ rbzero.trace_state\[2\] vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__buf_4
XFILLER_136_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18830_ rbzero.pov.spi_buffer\[24\] rbzero.pov.ready_buffer\[24\] _02989_ vssd1 vssd1
+ vccd1 vccd1 _02995_ sky130_fd_sc_hd__mux2_1
X_11165_ _04214_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15973_ _09024_ _09067_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__xnor2_1
X_11096_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _04340_ vssd1 vssd1 vccd1 vccd1 _04348_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18761_ _02952_ _02954_ _02955_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__nor3_1
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17712_ _10059_ _09243_ _01776_ _01887_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__o31a_1
X_14924_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.trackDistX\[-2\] _08062_
+ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__mux2_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _02889_ _02890_ _02860_ _02864_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o2111a_1
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _01931_ _01932_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__and2_1
X_14855_ _06470_ _08009_ _08010_ _07891_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__a31o_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _06936_ _06974_ _06976_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__a21bo_1
X_17574_ _01754_ _01756_ _01865_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a21boi_2
XFILLER_205_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14786_ _06580_ _07815_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__or2_1
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ rbzero.tex_r1\[13\] _05185_ _05186_ _04937_ vssd1 vssd1 vccd1 vccd1 _05187_
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ _09005_ _09242_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__nor2_1
X_19313_ rbzero.spi_registers.new_texadd\[3\]\[23\] _03239_ _03270_ _03265_ vssd1
+ vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__o211a_1
XFILLER_182_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13737_ _06889_ _06899_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__xnor2_1
X_10949_ _04271_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16456_ _08516_ _09037_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__nor2_1
X_19244_ rbzero.spi_registers.new_texadd\[2\]\[17\] _03221_ _03231_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__o211a_1
X_13668_ _06835_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__xor2_1
XFILLER_32_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15407_ _08039_ _08161_ _08398_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__or3_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ net20 net21 vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__and2b_1
X_19175_ rbzero.spi_registers.texadd1\[12\] _03189_ vssd1 vssd1 vccd1 vccd1 _03192_
+ sky130_fd_sc_hd__or2_1
X_16387_ _09340_ _09342_ _09465_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__a21oi_1
X_13599_ _06754_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__nor2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18126_ _02394_ _02396_ _02395_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a21boi_1
X_15338_ _08430_ _08432_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__nand2_1
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__or2_1
X_15269_ _08355_ _08361_ _08363_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__o21ai_1
X_17008_ _10027_ _10028_ vssd1 vssd1 vccd1 vccd1 _10029_ sky130_fd_sc_hd__nand2_1
XFILLER_160_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18959_ rbzero.spi_registers.spi_buffer\[10\] rbzero.spi_registers.spi_buffer\[9\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21970_ net496 _01559_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20921_ clknet_leaf_52_i_clk _00510_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20852_ clknet_leaf_50_i_clk _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20783_ _03110_ _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__and3_1
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21404_ clknet_leaf_32_i_clk _00993_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21335_ clknet_leaf_31_i_clk _00924_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_leak
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19695__73 clknet_1_0__leaf__03462_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XFILLER_190_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21266_ clknet_leaf_27_i_clk _00855_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20217_ _03775_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
X_21197_ clknet_leaf_29_i_clk _00786_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20148_ _05644_ _03734_ _03726_ _03736_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a22o_1
XFILLER_131_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20079_ _05120_ _03685_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__or2_1
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ rbzero.map_overlay.i_mapdx\[0\] _06144_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nor2_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03804_ clknet_0__03804_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03804_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _05093_ _05100_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__and2b_2
XFILLER_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _06613_ _07808_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__o21ba_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ rbzero.row_render.wall\[1\] rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1
+ vccd1 _05042_ sky130_fd_sc_hd__and2b_1
XFILLER_61_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _04194_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__clkbuf_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14571_ _07717_ _07739_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__o21bai_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _04913_ vssd1 vssd1 vccd1 vccd1 _04973_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16310_ _09400_ _09401_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__nor2_1
XFILLER_202_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _06687_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nor2_2
XFILLER_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17290_ _10188_ _10197_ _10196_ vssd1 vssd1 vccd1 vccd1 _10309_ sky130_fd_sc_hd__a21o_1
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _04158_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _09143_ _09216_ _09214_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13453_ _06451_ _06455_ _06603_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10665_ rbzero.tex_r0\[4\] rbzero.tex_r0\[3\] _04121_ vssd1 vssd1 vccd1 vccd1 _04122_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _05198_ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__or2_1
XFILLER_167_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16172_ _09241_ _09264_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__xor2_1
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13384_ _06439_ _06440_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__nor2_1
X_10596_ _04085_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15123_ _08185_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__buf_4
X_12335_ _04946_ _05518_ _05519_ _05520_ _04890_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__o221a_1
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15054_ _06260_ vssd1 vssd1 vccd1 vccd1 _08149_ sky130_fd_sc_hd__buf_6
X_19931_ rbzero.debug_overlay.playerX\[0\] _03559_ _03590_ _03584_ vssd1 vssd1 vccd1
+ vccd1 _01176_ sky130_fd_sc_hd__a211o_1
X_12266_ rbzero.tex_g1\[32\] _04934_ _04932_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_
+ sky130_fd_sc_hd__a31o_1
XFILLER_135_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14005_ _07174_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__nand2_1
X_11217_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__inv_2
X_19862_ _03543_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__buf_2
X_12197_ rbzero.tex_g1\[14\] _05236_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__or2_1
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03462_ _03462_ vssd1 vssd1 vccd1 vccd1 clknet_0__03462_ sky130_fd_sc_hd__clkbuf_16
X_18813_ rbzero.pov.spi_buffer\[16\] rbzero.pov.ready_buffer\[16\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11148_ _04375_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__clkbuf_1
X_19793_ _03507_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18744_ rbzero.spi_registers.spi_counter\[2\] rbzero.spi_registers.spi_counter\[1\]
+ _02936_ _02931_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__or4_1
XFILLER_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _04259_ vssd1 vssd1 vccd1 vccd1 _04339_
+ sky130_fd_sc_hd__mux2_1
X_15956_ _08148_ _09049_ _09050_ _08454_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__a31o_1
XFILLER_209_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14907_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.trackDistX\[-7\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__mux2_1
X_15887_ _08976_ _08980_ _08981_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__or3_1
XFILLER_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18675_ _02821_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02876_
+ sky130_fd_sc_hd__xnor2_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17626_ _01915_ _01916_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14838_ rbzero.wall_tracer.stepDistY\[1\] _07996_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _07997_ sky130_fd_sc_hd__mux2_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _01734_ _01736_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__nor2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14769_ rbzero.wall_tracer.stepDistY\[-7\] _07935_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07936_ sky130_fd_sc_hd__mux2_1
XFILLER_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _09477_ _09598_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__xnor2_1
X_17488_ _01778_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__xnor2_1
X_20539__381 clknet_1_1__leaf__03806_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__inv_2
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19227_ _03207_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__buf_2
X_16439_ _08813_ _08497_ _08409_ _09528_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__o22a_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19158_ rbzero.spi_registers.texadd1\[5\] _03176_ vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__or2_1
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__nand2_1
XFILLER_172_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19089_ rbzero.spi_registers.got_new_texadd\[0\] _03100_ vssd1 vssd1 vccd1 vccd1
+ _03142_ sky130_fd_sc_hd__and2_1
XFILLER_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21120_ clknet_leaf_91_i_clk _00709_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21051_ clknet_leaf_95_i_clk _00640_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20002_ _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__inv_2
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20284__151 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__inv_2
XFILLER_28_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21953_ net479 _01542_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ clknet_leaf_41_i_clk _00493_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21884_ net410 _01473_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20835_ clknet_leaf_66_i_clk _00424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20766_ _02749_ _02748_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__nor2_1
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20697_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03913_
+ sky130_fd_sc_hd__or2_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10450_ rbzero.tex_r1\[39\] net73 _04002_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ rbzero.tex_g0\[2\] _05195_ _05185_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a21o_1
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21318_ clknet_leaf_30_i_clk _00907_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12051_ rbzero.tex_r1\[35\] _04924_ _05239_ _04944_ vssd1 vssd1 vccd1 vccd1 _05240_
+ sky130_fd_sc_hd__o211a_1
X_21249_ clknet_leaf_26_i_clk _00838_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20367__226 clknet_1_1__leaf__03789_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__inv_2
XFILLER_172_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11002_ rbzero.tex_b1\[35\] rbzero.tex_b1\[36\] _04292_ vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15810_ _08865_ _08904_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__xnor2_1
X_16790_ _09818_ _09819_ _09817_ vssd1 vssd1 vccd1 vccd1 _09821_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _08796_ _08798_ _08797_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__a21o_1
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__clkinv_2
XFILLER_133_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11904_ _05076_ _05088_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a21o_4
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15672_ _08195_ _08250_ _08251_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__or3b_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _02534_ _02685_ _02686_ _09745_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a31o_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _06010_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nand2_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _01702_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__xor2_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _07625_ _07673_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__nor2_1
X_11835_ _04812_ _04917_ _04826_ _05024_ _05021_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__a32o_1
X_18391_ _02621_ _02622_ rbzero.wall_tracer.rayAddendX\[3\] _09744_ vssd1 vssd1 vccd1
+ vccd1 _02623_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _10271_ _10360_ vssd1 vssd1 vccd1 vccd1 _10361_ sky130_fd_sc_hd__nand2_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14554_ _07689_ _07724_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__xor2_1
XFILLER_18_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _04941_ _04945_ _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a211o_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _06604_ _06608_ _06554_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__mux2_1
XFILLER_105_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17273_ _08580_ _08382_ _08617_ _09076_ vssd1 vssd1 vccd1 vccd1 _10292_ sky130_fd_sc_hd__or4_1
XFILLER_158_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10717_ _04149_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__clkbuf_1
X_14485_ _06729_ _07310_ _07655_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__a21o_1
X_11697_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__buf_6
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ _08733_ _09314_ _09316_ _09193_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__a31o_1
X_19012_ _04687_ _05651_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__and3_1
X_13436_ _06463_ _06465_ _06603_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__mux2_1
X_10648_ rbzero.tex_r0\[12\] rbzero.tex_r0\[11\] _04110_ vssd1 vssd1 vccd1 vccd1 _04113_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19659__40 clknet_1_0__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ _08335_ _09076_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__nor2_1
X_13367_ _06516_ _06526_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__nor2_1
X_10579_ _04076_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ rbzero.wall_tracer.stepDistX\[-4\] _06262_ _08200_ vssd1 vssd1 vccd1 vccd1
+ _08201_ sky130_fd_sc_hd__o21bai_4
X_12318_ _04952_ _05499_ _05503_ _04889_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a211o_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16086_ _09178_ _09179_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__xnor2_1
X_13298_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__buf_4
X_19674__54 clknet_1_1__leaf__03460_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15037_ _04432_ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__buf_4
X_19914_ _08279_ _03570_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__nor2_1
X_12249_ _05429_ _05431_ _05433_ _05435_ _04812_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__o221a_1
XFILLER_130_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19845_ rbzero.pov.spi_buffer\[59\] rbzero.pov.spi_buffer\[60\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03535_ sky130_fd_sc_hd__mux2_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19776_ _03498_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16988_ _10006_ _10009_ vssd1 vssd1 vccd1 vccd1 _10010_ sky130_fd_sc_hd__xnor2_4
X_18727_ _02922_ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15939_ _09025_ _09032_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__or2_1
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18658_ _05127_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02860_
+ sky130_fd_sc_hd__nand2_1
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17609_ rbzero.wall_tracer.visualWallDist\[4\] _08421_ _01699_ _01899_ vssd1 vssd1
+ vccd1 vccd1 _01900_ sky130_fd_sc_hd__a31o_1
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18589_ _02794_ rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02796_
+ sky130_fd_sc_hd__and2_1
XFILLER_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20620_ _03734_ _03847_ _03848_ _03740_ rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1
+ _01607_ sky130_fd_sc_hd__a32o_1
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__05879_ _05879_ vssd1 vssd1 vccd1 vccd1 clknet_0__05879_ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21103_ clknet_leaf_72_i_clk _00692_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21034_ clknet_leaf_46_i_clk _00623_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21936_ net462 _01525_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21867_ net393 _01456_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11620_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__buf_8
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20818_ clknet_leaf_63_i_clk _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21798_ net324 _01387_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ _04733_ _04734_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and3_1
X_20749_ _03728_ _03938_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__and3_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10502_ rbzero.tex_r1\[14\] rbzero.tex_r1\[15\] _04024_ vssd1 vssd1 vccd1 vccd1 _04034_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14270_ _07419_ _07427_ _07440_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__inv_2
XFILLER_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ _06359_ _06361_ _06365_ _06386_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__a2111o_2
X_10433_ rbzero.tex_r1\[47\] rbzero.tex_r1\[48\] _03991_ vssd1 vssd1 vccd1 vccd1 _03998_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__inv_2
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12103_ _04722_ _04729_ _04719_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__o21bai_1
XFILLER_174_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17960_ _02152_ _02246_ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a21o_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ rbzero.trace_state\[3\] rbzero.trace_state\[2\] vssd1 vssd1 vccd1 vccd1 _06259_
+ sky130_fd_sc_hd__and2b_1
XFILLER_3_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16911_ _08151_ _08580_ vssd1 vssd1 vccd1 vccd1 _09933_ sky130_fd_sc_hd__nor2_1
X_12034_ rbzero.tex_r1\[24\] _05185_ _05181_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_
+ sky130_fd_sc_hd__a31o_1
XFILLER_105_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17891_ _01984_ _01987_ _01985_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__o21a_1
XFILLER_137_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19630_ rbzero.pov.spi_counter\[2\] _03442_ _03440_ vssd1 vssd1 vccd1 vccd1 _03449_
+ sky130_fd_sc_hd__o21ai_1
X_16842_ _09863_ _09864_ _09866_ vssd1 vssd1 vccd1 vccd1 _09867_ sky130_fd_sc_hd__a21o_1
XFILLER_19_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19561_ rbzero.spi_registers.new_texadd\[0\]\[22\] rbzero.spi_registers.spi_buffer\[22\]
+ _03380_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
X_16773_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ _09805_ vssd1 vssd1 vccd1 vccd1 _09806_ sky130_fd_sc_hd__a21o_1
X_13985_ _07055_ _07057_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18512_ _06117_ _09785_ _02728_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15724_ _08766_ _08817_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__xor2_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ rbzero.debug_overlay.playerY\[2\] vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__inv_2
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19492_ rbzero.spi_registers.new_mapd\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _03361_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _02597_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _02671_
+ sky130_fd_sc_hd__and2_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20421__275 clknet_1_0__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__inv_2
X_15655_ _08726_ _08749_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__nor2_1
X_12867_ _06018_ _06024_ _06028_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a21oi_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _05006_ _05007_ _04944_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__mux2_1
XFILLER_178_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14606_ _07770_ _07775_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__or2_1
X_15586_ _08245_ _08275_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__nor2_1
X_18374_ _08136_ _02605_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a21o_1
X_12798_ _05952_ _05966_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__a21o_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _10342_ _10343_ vssd1 vssd1 vccd1 vccd1 _10344_ sky130_fd_sc_hd__xnor2_1
X_14537_ _07683_ _07706_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__nor2_1
XFILLER_105_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ _04814_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__clkbuf_8
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17256_ _09520_ _09362_ vssd1 vssd1 vccd1 vccd1 _10275_ sky130_fd_sc_hd__nor2_1
X_14468_ _06993_ _07476_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__or2_1
XFILLER_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16207_ _09298_ _09299_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__and2_1
XFILLER_146_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13419_ _06571_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__clkbuf_4
X_17187_ _08816_ _09560_ _10082_ vssd1 vssd1 vccd1 vccd1 _10207_ sky130_fd_sc_hd__or3b_1
X_14399_ _07556_ _07567_ _07569_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__a21oi_1
X_16138_ _09229_ _09231_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__or2_1
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _09145_ _09033_ _09161_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__nand3_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19828_ rbzero.pov.spi_buffer\[51\] rbzero.pov.spi_buffer\[52\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XFILLER_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19759_ _03489_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21721_ net247 _01310_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20396__252 clknet_1_0__leaf__03792_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__inv_2
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21652_ clknet_leaf_96_i_clk _01241_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20603_ _03734_ _03833_ _03834_ _03814_ rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1
+ _01604_ sky130_fd_sc_hd__a32o_1
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21583_ clknet_leaf_91_i_clk _01172_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20534_ clknet_1_0__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__buf_1
XFILLER_123_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_79 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_79/HI o_rgb[4] sky130_fd_sc_hd__conb_1
XFILLER_181_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19653__35 clknet_1_0__leaf__03458_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
XFILLER_134_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22066_ clknet_leaf_36_i_clk _01655_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21017_ clknet_leaf_74_i_clk _00606_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_43_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20566__26 clknet_1_0__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
X_13770_ _06728_ _06737_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__nor2_1
X_10982_ _04288_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_40_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12721_ net29 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__inv_2
X_21919_ net445 _01508_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15440_ _08340_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_2_0_0_i_clk clknet_1_0_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12652_ net23 _05829_ net25 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a21o_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _04762_ _04766_ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__o21bai_4
XFILLER_12_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15371_ _08462_ _08465_ _08357_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__a21o_2
XFILLER_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12583_ net16 vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_168_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17110_ _10128_ _10129_ _10130_ vssd1 vssd1 vccd1 vccd1 _10131_ sky130_fd_sc_hd__and3_1
X_14322_ _07432_ _07489_ _07492_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__o21ai_1
X_11534_ rbzero.map_overlay.i_mapdx\[0\] _04413_ _04414_ rbzero.map_overlay.i_mapdx\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a22o_1
X_18090_ _02369_ _02370_ _02364_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__o21a_1
XFILLER_129_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _10060_ _10061_ vssd1 vssd1 vccd1 vccd1 _10062_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14253_ _07417_ _07366_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__or2_1
X_11465_ _04651_ _04652_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__nand2_1
XFILLER_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _06299_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__and2_1
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10416_ rbzero.tex_r1\[55\] rbzero.tex_r1\[56\] _03980_ vssd1 vssd1 vccd1 vccd1 _03989_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14184_ _07343_ _07354_ _07352_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11396_ _04575_ _04521_ _04585_ _04587_ _03971_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__o311a_1
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13135_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__nor2_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _02475_ _02474_ _03078_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_152_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17943_ _02229_ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__xnor2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ rbzero.map_overlay.i_otherx\[3\] _06228_ vssd1 vssd1 vccd1 vccd1 _06242_
+ sky130_fd_sc_hd__nor2_1
XFILLER_112_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _05197_ _05201_ _05203_ _05205_ _04955_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__o221a_1
XFILLER_94_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17874_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__nand2_1
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19613_ _03435_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__clkbuf_1
X_16825_ _06104_ _09227_ vssd1 vssd1 vccd1 vccd1 _09852_ sky130_fd_sc_hd__nand2_1
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19544_ _03400_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16756_ rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\] _09118_ vssd1 vssd1
+ vccd1 vccd1 _09792_ sky130_fd_sc_hd__o21a_1
XFILLER_207_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13968_ _07081_ _07131_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__o21a_1
XFILLER_185_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15707_ _08773_ _08778_ _08781_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__and3_1
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _06086_ _06087_ _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__o21ai_1
X_19475_ _03364_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13899_ _06942_ _06722_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__nor2_1
X_16687_ rbzero.row_render.size\[10\] _09752_ _09754_ _08000_ vssd1 vssd1 vccd1 vccd1
+ _00493_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ _02653_ _02654_ _02642_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a21o_1
X_15638_ rbzero.wall_tracer.visualWallDist\[-9\] _08149_ _08357_ rbzero.debug_overlay.playerX\[-9\]
+ _08438_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__a221o_4
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18357_ _02574_ _02590_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15569_ _08178_ _08440_ _08636_ _08638_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17308_ _10311_ _10326_ vssd1 vssd1 vccd1 vccd1 _10327_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18288_ _02525_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__buf_4
XFILLER_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17239_ _09822_ _10258_ vssd1 vssd1 vccd1 vccd1 _10259_ sky130_fd_sc_hd__nand2_1
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20181_ rbzero.spi_registers.new_texadd\[3\]\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21704_ net230 _01293_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21635_ clknet_leaf_82_i_clk _01224_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21566_ clknet_leaf_94_i_clk _01155_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21497_ clknet_leaf_97_i_clk _01086_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11181_ _04392_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20379_ clknet_1_0__leaf__03785_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__buf_1
XFILLER_162_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22049_ clknet_leaf_39_i_clk _01638_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14940_ _08065_ _08073_ _08074_ _08061_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__o211a_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14871_ rbzero.wall_tracer.stepDistY\[7\] _08023_ _07983_ vssd1 vssd1 vccd1 vccd1
+ _08024_ sky130_fd_sc_hd__mux2_1
XFILLER_29_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16610_ _09697_ _09699_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _06755_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__clkbuf_4
X_17590_ _01784_ _01799_ _01797_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a21o_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16541_ _09499_ _09630_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__xor2_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13753_ _06914_ _06922_ _06923_ _06849_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__o211a_1
X_10965_ _04279_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12704_ _05881_ _05057_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__or2_1
X_19260_ rbzero.spi_registers.got_new_texadd\[3\] _03100_ vssd1 vssd1 vccd1 vccd1
+ _03241_ sky130_fd_sc_hd__and2_1
XFILLER_188_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13684_ _06854_ _06721_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__nand2_1
X_16472_ _08011_ _08023_ _08449_ _09188_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__or4_1
X_10896_ _04243_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18211_ rbzero.spi_registers.spi_cmd\[2\] vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__clkbuf_2
X_15423_ _08253_ _08373_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__nor2_1
X_12635_ net44 _05791_ _05790_ _05808_ _05053_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__a32o_1
X_19191_ rbzero.spi_registers.new_texadd\[1\]\[19\] _03188_ _03200_ _03197_ vssd1
+ vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__o211a_1
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03800_ clknet_0__03800_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03800_
+ sky130_fd_sc_hd__clkbuf_16
X_18142_ _02341_ _02414_ _02415_ _02339_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__o31a_1
X_15354_ _07992_ _08393_ _08006_ _08000_ _07996_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__a2111o_1
XFILLER_180_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12566_ _05726_ _05745_ _05721_ _05746_ net14 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a221o_1
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14305_ _07158_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__clkbuf_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11517_ rbzero.map_overlay.i_otherx\[3\] _04410_ _04704_ _04705_ _04706_ vssd1 vssd1
+ vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
XFILLER_102_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20533__376 clknet_1_0__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__inv_2
X_18073_ _02353_ _02354_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__and3_1
X_15285_ _07975_ _08147_ _08379_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__a21oi_2
X_12497_ _04589_ _04704_ _04419_ _03973_ _05646_ net5 vssd1 vssd1 vccd1 vccd1 _05679_
+ sky130_fd_sc_hd__mux4_1
XFILLER_176_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17024_ _10043_ _10044_ vssd1 vssd1 vccd1 vccd1 _10045_ sky130_fd_sc_hd__nand2_1
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14236_ _07404_ _07406_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__or2_1
X_20232__104 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__inv_2
X_11448_ gpout0.hpos\[4\] _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or2_2
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _07206_ _07310_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__or2b_1
X_11379_ _03971_ _04543_ _04570_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o21ai_1
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__nand2_1
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ rbzero.spi_registers.spi_buffer\[18\] rbzero.spi_registers.spi_buffer\[17\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
X_14098_ _07260_ _07222_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__and2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _02114_ _02097_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__or2b_1
XFILLER_6_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _06113_ _06224_ _06088_ _06144_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17857_ _02135_ _02145_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16808_ _09822_ _09105_ vssd1 vssd1 vccd1 vccd1 _09837_ sky130_fd_sc_hd__nand2_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17788_ _01965_ _01968_ _02076_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__and3_2
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19527_ _03391_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
X_16739_ _09764_ _09776_ vssd1 vssd1 vccd1 vccd1 _09777_ sky130_fd_sc_hd__and2_1
XFILLER_35_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19458_ rbzero.spi_registers.new_vshift\[3\] _02485_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03355_ sky130_fd_sc_hd__mux2_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18409_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _02598_
+ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o21ai_1
XFILLER_194_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19389_ _03315_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
X_21420_ clknet_leaf_4_i_clk _01009_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_175_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21351_ clknet_leaf_35_i_clk _00940_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21282_ clknet_leaf_100_i_clk _00871_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20164_ _03746_ _03744_ _03747_ _04409_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a211oi_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ rbzero.pov.ready_buffer\[21\] _03684_ _03701_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01229_ sky130_fd_sc_hd__o211a_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20328__190 clknet_1_1__leaf__03786_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__inv_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20997_ clknet_leaf_99_i_clk _00586_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ rbzero.tex_g1\[27\] rbzero.tex_g1\[28\] _04166_ vssd1 vssd1 vccd1 vccd1 _04167_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10681_ rbzero.tex_g1\[59\] rbzero.tex_g1\[60\] _04046_ vssd1 vssd1 vccd1 vccd1 _04130_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12420_ rbzero.tex_b1\[3\] _04927_ _04929_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__and3_1
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21618_ clknet_leaf_71_i_clk _01207_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12351_ _05531_ _05533_ _05536_ _04952_ _04889_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a221o_1
X_21549_ clknet_leaf_92_i_clk _01138_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ rbzero.spi_registers.texadd1\[6\] _04460_ _04469_ _04493_ vssd1 vssd1 vccd1
+ vccd1 _04494_ sky130_fd_sc_hd__a211o_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15070_ rbzero.wall_tracer.visualWallDist\[2\] _08149_ vssd1 vssd1 vccd1 vccd1 _08165_
+ sky130_fd_sc_hd__nand2_4
XFILLER_119_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12282_ _05176_ _05468_ _05051_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14021_ _07181_ _07191_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__or2_1
XFILLER_5_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__buf_2
XFILLER_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11164_ _04383_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18760_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ _02929_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and3_1
X_15972_ _09064_ _09066_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__xor2_1
X_11095_ _04347_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17711_ _01999_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__xor2_1
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14923_ _06217_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__clkbuf_4
X_18691_ _02862_ _02863_ _02876_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__or3_1
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17642_ _01931_ _01932_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__nor2_1
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _06631_ _07962_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__nand2_1
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13805_ _06729_ _06700_ _06808_ _06728_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__a22o_1
X_17573_ _01752_ _01753_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__or2_1
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11997_ _04831_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__buf_4
X_14785_ _07822_ _07811_ _07949_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__a21o_1
X_19312_ rbzero.spi_registers.texadd3\[23\] _03241_ vssd1 vssd1 vccd1 vccd1 _03270_
+ sky130_fd_sc_hd__or2_1
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16524_ _09008_ _09363_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__nor2_1
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10948_ rbzero.tex_b1\[61\] rbzero.tex_b1\[62\] _04270_ vssd1 vssd1 vccd1 vccd1 _04271_
+ sky130_fd_sc_hd__mux2_1
X_13736_ _06901_ _06903_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__a211o_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19243_ rbzero.spi_registers.texadd2\[17\] _03222_ vssd1 vssd1 vccd1 vccd1 _03231_
+ sky130_fd_sc_hd__or2_1
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ _09303_ _09545_ _09419_ _09416_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__a22o_1
X_10879_ _04234_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ _06836_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _08408_ _08440_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__nor2_1
XFILLER_129_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12618_ _05792_ _05765_ _05770_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__and3b_1
X_19174_ rbzero.spi_registers.new_texadd\[1\]\[11\] _03188_ _03191_ _03184_ vssd1
+ vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__o211a_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13598_ _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__clkbuf_4
X_16386_ _09472_ _09473_ _09470_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__o21ba_1
XFILLER_185_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18125_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__and2_1
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15337_ _08431_ _08429_ _08413_ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__o21bai_1
X_12549_ gpout0.vpos\[1\] net10 vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or2b_1
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18056_ _06104_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _08152_ _08171_ _08362_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__or3_2
XFILLER_67_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17007_ _09953_ _09930_ vssd1 vssd1 vccd1 vccd1 _10028_ sky130_fd_sc_hd__or2b_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14219_ _07380_ _07388_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__a21oi_1
X_15199_ _06065_ _06366_ rbzero.side_hot vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__mux2_1
XFILLER_126_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18958_ _03051_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__buf_4
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17909_ _08530_ _02105_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a21o_1
XFILLER_117_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18889_ rbzero.pov.spi_buffer\[52\] rbzero.pov.ready_buffer\[52\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
XFILLER_55_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20920_ clknet_leaf_53_i_clk _00509_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20851_ clknet_leaf_52_i_clk _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20782_ gpout2.clk_div\[1\] gpout2.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__or2_1
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20516__360 clknet_1_1__leaf__03804_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__inv_2
X_21403_ clknet_leaf_27_i_clk _00992_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21334_ clknet_leaf_31_i_clk _00923_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21265_ clknet_leaf_25_i_clk _00854_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20216_ rbzero.spi_registers.new_texadd\[3\]\[23\] rbzero.spi_registers.spi_buffer\[23\]
+ _03384_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__mux2_1
XFILLER_173_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21196_ clknet_leaf_29_i_clk _00785_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20147_ _05644_ _03092_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__o21a_1
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03803_ clknet_0__03803_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03803_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ rbzero.pov.ready_buffer\[13\] _03684_ _03692_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01221_ sky130_fd_sc_hd__o211a_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11920_ _05106_ _05107_ _05108_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1
+ vccd1 _05109_ sky130_fd_sc_hd__a22o_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20261__130 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__inv_2
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _05020_ _05028_ _05030_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a31o_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ rbzero.tex_g1\[2\] rbzero.tex_g1\[3\] _04188_ vssd1 vssd1 vccd1 vccd1 _04194_
+ sky130_fd_sc_hd__mux2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _07640_ _07722_ _07740_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__nor3_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11782_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _04909_ vssd1 vssd1 vccd1 vccd1 _04972_
+ sky130_fd_sc_hd__mux2_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ rbzero.tex_g1\[35\] rbzero.tex_g1\[36\] _04155_ vssd1 vssd1 vccd1 vccd1 _04158_
+ sky130_fd_sc_hd__mux2_1
X_13521_ _06469_ _06689_ _06690_ _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__o31a_4
XFILLER_202_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _09267_ _09332_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__xnor2_1
X_13452_ _06619_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__and2_1
X_10664_ _04054_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__clkbuf_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12403_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _04893_ vssd1 vssd1 vccd1 vccd1 _05588_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16171_ _09244_ _09263_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__xnor2_1
X_13383_ _06540_ _06542_ _06545_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__nor4_4
X_10595_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _04077_ vssd1 vssd1 vccd1 vccd1 _04085_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12334_ rbzero.tex_b0\[19\] _04926_ _04928_ _05198_ vssd1 vssd1 vccd1 vccd1 _05520_
+ sky130_fd_sc_hd__a31o_1
X_15122_ _08215_ _08216_ vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__and2_1
XFILLER_86_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ rbzero.pov.ready_buffer\[68\] _03586_ _03588_ _03589_ _03569_ vssd1 vssd1
+ vccd1 vccd1 _03590_ sky130_fd_sc_hd__o221a_1
X_15053_ _08147_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__buf_4
X_12265_ rbzero.tex_g1\[33\] _04891_ _04830_ _04917_ vssd1 vssd1 vccd1 vccd1 _05452_
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ _07117_ _07173_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__nand2_1
X_11216_ gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19861_ rbzero.pov.spi_buffer\[67\] rbzero.pov.spi_buffer\[68\] _03534_ vssd1 vssd1
+ vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux2_1
X_12196_ _05383_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 o_gpout[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__buf_2
Xclkbuf_0__03461_ _03461_ vssd1 vssd1 vccd1 vccd1 clknet_0__03461_ sky130_fd_sc_hd__clkbuf_16
X_18812_ _02985_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
X_11147_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _04373_ vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__mux2_1
X_19792_ rbzero.pov.spi_buffer\[34\] rbzero.pov.spi_buffer\[35\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20344__205 clknet_1_0__leaf__03787_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__inv_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18743_ _02936_ _02931_ _02937_ _02938_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__o211ai_1
X_11078_ _04338_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
X_15955_ _08012_ _08450_ _08015_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__o21ai_1
XFILLER_3_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14906_ _08036_ _08049_ _08050_ _01633_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__o211a_1
XFILLER_209_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18674_ _09753_ _02865_ _02866_ _02875_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__a31o_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _08912_ _08943_ _08975_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _01882_ _01883_ _01914_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__nand3_1
X_14837_ _06669_ _07931_ _07995_ _06581_ _07866_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__o221ai_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ _01828_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
X_14768_ _07933_ _07934_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__nand2_2
XFILLER_108_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16507_ _09121_ _09597_ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__xor2_1
X_13719_ _06707_ _06807_ _06806_ _06809_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a22o_1
X_17487_ _09520_ _09491_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__nor2_1
XFILLER_177_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14699_ rbzero.wall_tracer.stepDistY\[-11\] _07867_ _07869_ vssd1 vssd1 vccd1 vccd1
+ _07870_ sky130_fd_sc_hd__mux2_1
X_19226_ _03205_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__clkbuf_4
X_16438_ _09528_ _08497_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__nor2_2
XFILLER_31_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19157_ rbzero.spi_registers.new_texadd\[1\]\[4\] _03174_ _03181_ _03169_ vssd1 vssd1
+ vccd1 vccd1 _00811_ sky130_fd_sc_hd__o211a_1
X_16369_ _09357_ _09460_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__xor2_1
XFILLER_157_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__nor2_1
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19088_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18039_ _02272_ _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__xnor2_1
X_21050_ clknet_leaf_87_i_clk _00639_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20001_ rbzero.debug_overlay.playerY\[3\] _03640_ _03436_ vssd1 vssd1 vccd1 vccd1
+ _03643_ sky130_fd_sc_hd__o21a_1
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21952_ net478 _01541_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ clknet_leaf_53_i_clk _00492_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21883_ net409 _01472_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20834_ clknet_leaf_66_i_clk _00423_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_165_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20765_ rbzero.wall_tracer.rayAddendY\[-9\] _09746_ _03950_ vssd1 vssd1 vccd1 vccd1
+ _01651_ sky130_fd_sc_hd__a21o_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20696_ _09732_ _03911_ _03912_ _03740_ rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1
+ _01619_ sky130_fd_sc_hd__a32o_1
XFILLER_126_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21317_ clknet_leaf_31_i_clk _00906_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ rbzero.tex_r1\[34\] _05236_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or2_1
X_21248_ clknet_leaf_25_i_clk _00837_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _04298_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21179_ clknet_leaf_13_i_clk _00768_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15740_ _08830_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__nor2_1
XFILLER_133_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ rbzero.debug_overlay.playerX\[5\] _06126_ rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\]
+ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a2111o_1
XFILLER_46_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11903_ _05076_ _05088_ _05069_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o21bai_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15671_ _08195_ _08275_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__or2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nand2_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _08499_ _08620_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14622_ _07713_ _07672_ _07790_ _07792_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__a22o_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\] vssd1 vssd1 vccd1
+ vccd1 _05024_ sky130_fd_sc_hd__nor2_1
X_18390_ _02618_ _02620_ _08135_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__o21ai_1
XFILLER_92_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _10358_ _10359_ vssd1 vssd1 vccd1 vccd1 _10360_ sky130_fd_sc_hd__xor2_1
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _04889_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__buf_4
XFILLER_144_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14553_ _07701_ _07700_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__nand2_1
XFILLER_199_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10716_ rbzero.tex_g1\[43\] rbzero.tex_g1\[44\] _04144_ vssd1 vssd1 vccd1 vccd1 _04149_
+ sky130_fd_sc_hd__mux2_1
X_13504_ _06641_ _06672_ _06674_ _06669_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__a211o_1
X_17272_ _08580_ _08618_ _09079_ _08382_ vssd1 vssd1 vccd1 vccd1 _10291_ sky130_fd_sc_hd__o22ai_1
XFILLER_202_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11696_ _04806_ _04822_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__or2_4
X_14484_ _07423_ _07248_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nor2_1
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19011_ _05653_ _05652_ _04642_ _05645_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__and4b_2
X_16223_ _08581_ _09315_ _09195_ _08461_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__o22ai_1
XFILLER_146_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10647_ _04112_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _06604_ _06605_ _06576_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__mux2_1
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16154_ _09246_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__inv_2
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ _06494_ _06527_ _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or3_4
X_10578_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _04066_ vssd1 vssd1 vccd1 vccd1 _04076_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ rbzero.wall_tracer.stepDistY\[-4\] _08157_ _08196_ _08199_ vssd1 vssd1 vccd1
+ vccd1 _08200_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12317_ _04826_ _05500_ _05501_ _05502_ _04939_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__o221a_1
XFILLER_127_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16085_ _09044_ _09046_ _08390_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13297_ _06448_ _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__and2_1
XFILLER_114_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ rbzero.tex_g1\[56\] _04934_ _04932_ _05434_ vssd1 vssd1 vccd1 vccd1 _05435_
+ sky130_fd_sc_hd__a31o_1
X_19913_ rbzero.debug_overlay.playerX\[-4\] _03569_ _03576_ _03302_ vssd1 vssd1 vccd1
+ vccd1 _01172_ sky130_fd_sc_hd__o211a_1
XFILLER_64_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15036_ _08132_ rbzero.mapdxw\[1\] _06151_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__mux2_1
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19844_ _03466_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__buf_4
X_12179_ _05364_ _05365_ _05366_ _05191_ _04953_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__o221a_1
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19775_ rbzero.pov.spi_buffer\[26\] rbzero.pov.spi_buffer\[27\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
XFILLER_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16987_ _09479_ _09592_ _10007_ _10008_ vssd1 vssd1 vccd1 vccd1 _10009_ sky130_fd_sc_hd__o31a_4
XFILLER_111_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18726_ _02822_ rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 _02923_
+ sky130_fd_sc_hd__xnor2_1
X_15938_ _09025_ _09032_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__nand2_1
XFILLER_110_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18657_ _02859_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15869_ _08431_ _08344_ _08696_ _08910_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__o22a_1
XFILLER_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17608_ _08428_ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__nor2_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18588_ _02794_ rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__nor2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17539_ _09167_ _10342_ _10331_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__o21ai_4
XFILLER_205_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19209_ _08116_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__buf_6
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21102_ clknet_leaf_71_i_clk _00691_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21033_ clknet_leaf_46_i_clk _00622_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21935_ net461 _01524_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ net392 _01455_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ clknet_leaf_60_i_clk _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21797_ net323 _01386_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11550_ _04735_ rbzero.map_overlay.i_mapdy\[0\] _04737_ rbzero.map_overlay.i_mapdy\[4\]
+ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o221a_1
XFILLER_184_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20748_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or2_1
XFILLER_156_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ _04033_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__clkbuf_1
X_20373__231 clknet_1_0__leaf__03790_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__inv_2
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ rbzero.debug_overlay.playerX\[1\] vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__inv_2
X_20679_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03898_
+ sky130_fd_sc_hd__or2_1
XFILLER_11_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13220_ _06389_ _06390_ _06323_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__mux2_2
X_10432_ _03997_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _06284_ _06320_ _04443_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__o211a_4
XFILLER_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _04744_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__and2_1
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _06217_ _06257_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and2b_1
XFILLER_105_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16910_ _09664_ _09675_ _09931_ vssd1 vssd1 vccd1 vccd1 _09932_ sky130_fd_sc_hd__a21bo_1
X_12033_ rbzero.tex_r1\[25\] _04982_ _05032_ _04919_ vssd1 vssd1 vccd1 vccd1 _05222_
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17890_ _02177_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__nand2_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _06103_ vssd1 vssd1 vccd1 vccd1 _09866_ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19560_ _03408_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__clkbuf_1
X_16772_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ _08123_ vssd1 vssd1 vccd1 vccd1 _09805_ sky130_fd_sc_hd__o21ai_1
X_13984_ _07058_ _07106_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__xor2_1
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18511_ _04671_ _08124_ _09844_ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__o211a_1
X_15723_ _08228_ _08336_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__or2_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19491_ _03372_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
X_12935_ rbzero.debug_overlay.playerY\[1\] vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__inv_2
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18442_ _02597_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _02670_
+ sky130_fd_sc_hd__nor2_1
X_15654_ _08716_ _08723_ _08725_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__and3_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12866_ _06026_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__inv_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20456__306 clknet_1_0__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__inv_2
X_14605_ _07770_ _07775_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__nand2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _04909_ vssd1 vssd1 vccd1 vccd1 _05007_
+ sky130_fd_sc_hd__mux2_1
X_18373_ _09744_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__buf_6
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15585_ _08663_ _08679_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__xor2_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ net38 _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nand2_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17324_ _09167_ _10330_ vssd1 vssd1 vccd1 vccd1 _10343_ sky130_fd_sc_hd__nor2_1
XFILLER_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14536_ _07683_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nand2_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _04923_ _04925_ _04930_ _04936_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__o221a_1
XFILLER_144_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17255_ _10180_ _10200_ _10273_ vssd1 vssd1 vccd1 vccd1 _10274_ sky130_fd_sc_hd__a21bo_1
XFILLER_159_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14467_ _07636_ _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__nand2_1
X_11679_ rbzero.row_render.size\[1\] _04449_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__and2_1
X_16206_ _09177_ _09180_ _09297_ _09292_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__a211o_1
X_13418_ _06554_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17186_ _09681_ _10204_ _10205_ _10088_ vssd1 vssd1 vccd1 vccd1 _10206_ sky130_fd_sc_hd__o22a_1
XFILLER_190_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14398_ _07564_ _07568_ _07566_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _09104_ _09116_ _09230_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13349_ _06477_ _06482_ _06489_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__or4_2
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16068_ _09145_ _09033_ _09161_ vssd1 vssd1 vccd1 vccd1 _09162_ sky130_fd_sc_hd__a21o_1
XFILLER_170_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15019_ _08117_ _05470_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__and2_1
XFILLER_155_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19827_ _03525_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19758_ rbzero.pov.spi_buffer\[18\] rbzero.pov.spi_buffer\[19\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18709_ _02794_ rbzero.debug_overlay.vplaneY\[-1\] _02822_ vssd1 vssd1 vccd1 vccd1
+ _02908_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21720_ net246 _01309_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21651_ clknet_leaf_85_i_clk _01240_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20602_ _03830_ _03831_ _03832_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__or3_1
XFILLER_178_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21582_ clknet_leaf_91_i_clk _01171_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_178_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22065_ clknet_leaf_79_i_clk _01654_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21016_ clknet_3_5_0_i_clk _00605_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10981_ rbzero.tex_b1\[45\] rbzero.tex_b1\[46\] _04281_ vssd1 vssd1 vccd1 vccd1 _04288_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12720_ net33 _05892_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and3_1
X_21918_ net444 _01507_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12651_ net27 _05828_ net23 _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and4b_1
XFILLER_43_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21849_ net375 _01438_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ _04767_ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__nor2_1
XFILLER_130_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12582_ _05762_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15370_ _08148_ _08463_ _08464_ _08454_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__a31o_1
XFILLER_141_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _06993_ _07204_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__o21bai_1
X_11533_ rbzero.map_overlay.i_mapdx\[2\] _04704_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__xor2_1
XFILLER_156_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _08151_ _08399_ vssd1 vssd1 vccd1 vccd1 _10061_ sky130_fd_sc_hd__nor2_2
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ _06792_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__clkbuf_4
X_11464_ _04651_ _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__or2_1
XFILLER_183_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _03988_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__clkbuf_1
X_13203_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__or2_1
XFILLER_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11395_ _04449_ _04513_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__or3_1
X_14183_ _07352_ _07353_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nor2_1
XFILLER_124_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13134_ _06297_ _06298_ _06303_ _06304_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__o31ai_4
XFILLER_139_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18991_ _03080_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17942_ _09662_ _02012_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__nor2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ rbzero.map_overlay.i_otherx\[4\] _06129_ _06089_ rbzero.map_overlay.i_othery\[1\]
+ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__a221o_1
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ rbzero.tex_r1\[0\] _05185_ _05181_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17873_ _02090_ _02160_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__or2_1
XFILLER_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19612_ rbzero.spi_registers.new_texadd\[1\]\[23\] rbzero.spi_registers.spi_buffer\[23\]
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
X_16824_ _09849_ _09850_ vssd1 vssd1 vccd1 vccd1 _09851_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19543_ rbzero.spi_registers.new_texadd\[0\]\[13\] rbzero.spi_registers.spi_buffer\[13\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _09778_ _09777_ _09787_ vssd1 vssd1 vccd1 vccd1 _09791_ sky130_fd_sc_hd__and3_1
XFILLER_4_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13967_ _07091_ _07137_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15706_ _08746_ _08784_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__a21o_1
XFILLER_98_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12918_ _06092_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__nand2_1
X_19474_ rbzero.spi_registers.new_mapd\[1\] _02481_ _03362_ vssd1 vssd1 vccd1 vccd1
+ _03364_ sky130_fd_sc_hd__mux2_1
XFILLER_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16686_ rbzero.row_render.size\[9\] _09752_ _09754_ _07996_ vssd1 vssd1 vccd1 vccd1
+ _00492_ sky130_fd_sc_hd__a22o_1
X_13898_ _06741_ _07066_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__a21oi_2
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18425_ _02597_ _05106_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__nand2_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15637_ _08229_ _08731_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__nor2_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _05997_ _05996_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__nand2_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18356_ _02588_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__nor2_1
X_15568_ _08641_ _08643_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__xnor2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17307_ _10317_ _10325_ vssd1 vssd1 vccd1 vccd1 _10326_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14519_ _07657_ _07654_ _07656_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nand3_1
XFILLER_187_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18287_ _02526_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__clkbuf_1
X_15499_ _08585_ _08507_ _08587_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__a21bo_1
XFILLER_163_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ _10254_ _10257_ vssd1 vssd1 vccd1 vccd1 _10258_ sky130_fd_sc_hd__and2_2
XFILLER_31_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17169_ _09044_ _09046_ _09528_ vssd1 vssd1 vccd1 vccd1 _10189_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20510__355 clknet_1_1__leaf__03803_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__inv_2
XFILLER_115_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20180_ _03756_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21703_ net229 _01292_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21634_ clknet_leaf_82_i_clk _01223_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21565_ clknet_leaf_92_i_clk _01154_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21496_ net214 _01085_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11180_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _04384_ vssd1 vssd1 vccd1 vccd1 _04392_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485__332 clknet_1_0__leaf__03801_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__inv_2
XFILLER_171_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22048_ clknet_leaf_39_i_clk _01637_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ _08021_ _08022_ _07891_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__a21o_1
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13821_ _06980_ _06989_ _06991_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__o21a_1
XFILLER_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16540_ _09627_ _09629_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__and2b_1
XFILLER_204_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _06846_ _06847_ _06848_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ rbzero.tex_b1\[53\] rbzero.tex_b1\[54\] _04270_ vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12703_ net28 vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__buf_2
X_16471_ _08471_ _09426_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__nand2_1
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13683_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__or2_2
XFILLER_44_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10895_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _04237_ vssd1 vssd1 vccd1 vccd1 _04243_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ rbzero.spi_registers.spi_cmd\[1\] vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__buf_2
X_15422_ _08370_ _08369_ _08516_ _08235_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__o22ai_1
X_12634_ net71 _05802_ _05803_ _05055_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a22o_1
X_19190_ rbzero.spi_registers.texadd1\[19\] _03189_ vssd1 vssd1 vccd1 vccd1 _03200_
+ sky130_fd_sc_hd__or2_1
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18141_ _02411_ _02412_ _02413_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15353_ _08441_ _08447_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__nor2_1
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _05053_ _05712_ _05715_ net44 vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a22o_1
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ _07460_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18072_ _02347_ _02348_ _02349_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__o21bai_1
X_11516_ gpout0.vpos\[4\] rbzero.map_overlay.i_othery\[1\] vssd1 vssd1 vccd1 vccd1
+ _04706_ sky130_fd_sc_hd__xor2_1
X_15284_ _08142_ _08378_ _08155_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__a21o_1
X_12496_ net7 _05640_ net8 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a21o_1
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ _08666_ _09079_ _09628_ vssd1 vssd1 vccd1 vccd1 _10044_ sky130_fd_sc_hd__or3_1
XFILLER_171_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _07327_ _07356_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ gpout0.hpos\[3\] _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__and2_1
XFILLER_171_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11378_ _04534_ _04540_ _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a21bo_1
X_14166_ _06720_ _07331_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__nor2_1
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__xor2_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18974_ _03071_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__clkbuf_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _06722_ _06640_ _06769_ _06720_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__or4_1
XFILLER_98_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17925_ _02134_ _02150_ _02148_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a21o_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _06157_ _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__nand2_1
XFILLER_121_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17856_ _02143_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__nor2_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _09834_ _09835_ vssd1 vssd1 vccd1 vccd1 _09836_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17787_ _01965_ _01968_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a21o_1
X_14999_ _08109_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ _09774_ _09775_ vssd1 vssd1 vccd1 vccd1 _09776_ sky130_fd_sc_hd__and2b_1
X_19526_ rbzero.spi_registers.new_texadd\[0\]\[5\] _02489_ _03381_ vssd1 vssd1 vccd1
+ vccd1 _03391_ sky130_fd_sc_hd__mux2_1
XFILLER_207_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19457_ _03354_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16669_ _04437_ _04433_ _05050_ _09747_ vssd1 vssd1 vccd1 vccd1 _09748_ sky130_fd_sc_hd__and4_1
XFILLER_167_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18408_ _02613_ _02625_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__or2b_1
XFILLER_72_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19388_ _02489_ rbzero.spi_registers.new_sky\[5\] _03309_ vssd1 vssd1 vccd1 vccd1
+ _03315_ sky130_fd_sc_hd__mux2_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18339_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__or2_1
XFILLER_33_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21350_ clknet_leaf_35_i_clk _00939_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20301_ clknet_1_1__leaf__03464_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__buf_1
XFILLER_162_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21281_ clknet_leaf_0_i_clk _00870_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20163_ _05652_ _04642_ _05645_ _03741_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__and4_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20094_ _02694_ _03655_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nand2_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20996_ clknet_leaf_1_i_clk _00585_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_69_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_168_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _04129_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21617_ clknet_leaf_71_i_clk _01206_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12350_ _05534_ _05535_ _04891_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__mux2_1
X_21548_ clknet_leaf_92_i_clk _01137_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ rbzero.spi_registers.texadd3\[6\] _04465_ _04455_ rbzero.spi_registers.texadd2\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a22o_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12281_ _04650_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__nor2_1
X_21479_ net197 _01068_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ _07182_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__xnor2_1
X_11232_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__buf_2
XFILLER_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _04373_ vssd1 vssd1 vccd1 vccd1 _04383_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15971_ _08419_ _08494_ _09065_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__a21boi_1
X_11094_ rbzero.tex_b0\[56\] rbzero.tex_b0\[55\] _04340_ vssd1 vssd1 vccd1 vccd1 _04347_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17710_ _09647_ _09621_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14922_ _08036_ _08059_ _08060_ _08061_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__o211a_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__inv_2
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _01818_ _09669_ _01817_ _01815_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o31a_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _06575_ _07986_ _08008_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__a21o_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _06936_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__nand2_1
X_17572_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__or2_1
X_14784_ _07822_ _07821_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__nor2_1
XFILLER_205_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11996_ _04982_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__buf_4
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19311_ rbzero.spi_registers.new_texadd\[3\]\[22\] _03239_ _03269_ _03265_ vssd1
+ vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__o211a_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16523_ _09540_ _09515_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__or2b_1
XFILLER_32_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ _06748_ _06761_ _06904_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__and3_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ _04143_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19242_ rbzero.spi_registers.new_texadd\[2\]\[16\] _03221_ _03230_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__o211a_1
X_16454_ _09053_ _09306_ _08910_ vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__a21oi_2
XFILLER_189_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13666_ _06722_ _06798_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__nor2_1
X_10878_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _04226_ vssd1 vssd1 vccd1 vccd1 _04234_
+ sky130_fd_sc_hd__mux2_1
X_15405_ _08499_ _08473_ _08458_ _08399_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__o22ai_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20550__11 clknet_1_1__leaf__03807_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
X_12617_ _05782_ _05789_ _05790_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a211o_1
X_19173_ rbzero.spi_registers.texadd1\[11\] _03189_ vssd1 vssd1 vccd1 vccd1 _03191_
+ sky130_fd_sc_hd__or2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ rbzero.texu_hot\[3\] _08145_ _09476_ _08085_ vssd1 vssd1 vccd1 vccd1 _00469_
+ sky130_fd_sc_hd__o211a_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _06710_ _06718_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__o21ai_1
XFILLER_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18124_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__nor2_1
X_15336_ _08390_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ _05703_ _05718_ _05723_ _05728_ _05707_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__o2111a_1
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _09804_ _02338_ _02340_ rbzero.wall_tracer.trackDistY\[-11\] vssd1 vssd1
+ vccd1 vccd1 _00550_ sky130_fd_sc_hd__o2bb2a_1
X_15267_ _08355_ _08361_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net7 vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__inv_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _09952_ _09932_ vssd1 vssd1 vccd1 vccd1 _10027_ sky130_fd_sc_hd__or2b_1
XFILLER_172_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14218_ _07383_ _07384_ _07387_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__and3_1
XFILLER_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15198_ _07919_ _07922_ _08143_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__a21o_1
XFILLER_141_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _07314_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__or2_1
XFILLER_28_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ _03062_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__clkbuf_1
X_17908_ _08814_ _09528_ _10093_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a21o_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18888_ _03025_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17839_ _10059_ _09621_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__nor2_1
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20850_ clknet_leaf_52_i_clk _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19509_ _02477_ _02930_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nor2_4
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20781_ gpout2.clk_div\[1\] gpout2.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__nand2_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21402_ clknet_leaf_27_i_clk _00991_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21333_ clknet_leaf_31_i_clk _00922_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21264_ clknet_leaf_25_i_clk _00853_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20215_ _03774_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21195_ clknet_leaf_29_i_clk _00784_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20146_ _05644_ _03092_ _04408_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20077_ rbzero.debug_overlay.vplaneX\[-7\] _03685_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__03802_ clknet_0__03802_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03802_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _05020_ _05039_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__nor2_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10801_ _04193_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__clkbuf_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _04969_ _04970_ _04944_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__mux2_1
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20979_ clknet_leaf_65_i_clk _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _06632_ _06631_ _06574_ _06628_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__or4_1
X_10732_ _04157_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13451_ _06620_ _06621_ _06554_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__mux2_1
X_10663_ _04120_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12402_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _05314_ vssd1 vssd1 vccd1 vccd1 _05587_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _09260_ _09262_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__xor2_1
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10594_ _04084_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__clkbuf_1
X_13382_ _06436_ _06548_ _06448_ _06549_ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a221o_1
XFILLER_16_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15121_ rbzero.debug_overlay.playerX\[-6\] _08207_ vssd1 vssd1 vccd1 vccd1 _08216_
+ sky130_fd_sc_hd__nand2_1
X_12333_ rbzero.tex_b0\[18\] _05314_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__and2_1
XFILLER_182_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15052_ _08146_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ rbzero.tex_g1\[35\] _04964_ _05450_ _04946_ vssd1 vssd1 vccd1 vccd1 _05451_
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _07117_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__or2_1
X_11215_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__buf_4
X_19860_ _03542_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
X_12195_ reg_rgb\[14\] _05382_ _05058_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_2
XFILLER_134_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_123_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__buf_2
Xclkbuf_0__03460_ _03460_ vssd1 vssd1 vccd1 vccd1 clknet_0__03460_ sky130_fd_sc_hd__clkbuf_16
X_18811_ rbzero.pov.spi_buffer\[15\] rbzero.pov.ready_buffer\[15\] _02978_ vssd1 vssd1
+ vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
XFILLER_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _04374_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__clkbuf_1
X_19791_ _03506_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11077_ net51 rbzero.tex_b0\[63\] _04259_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
X_18742_ rbzero.spi_registers.spi_counter\[2\] _02475_ rbzero.spi_registers.spi_cmd\[3\]
+ rbzero.spi_registers.spi_counter\[1\] vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__o31a_1
X_15954_ _08012_ _08015_ _08450_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__or3_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14905_ rbzero.wall_tracer.visualWallDist\[-8\] _08047_ vssd1 vssd1 vccd1 vccd1 _08050_
+ sky130_fd_sc_hd__or2_1
X_18673_ _02873_ _02874_ rbzero.wall_tracer.rayAddendY\[5\] _09744_ vssd1 vssd1 vccd1
+ vccd1 _02875_ sky130_fd_sc_hd__a2bb2o_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _08978_ _08979_ vssd1 vssd1 vccd1 vccd1 _08980_ sky130_fd_sc_hd__nor2_1
XFILLER_209_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _01882_ _01883_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a21o_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14836_ _06575_ _07862_ _07994_ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__o21ai_2
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17555_ _01845_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__nor2_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14767_ _06470_ _07826_ _07823_ _07891_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__a31oi_2
X_11979_ rbzero.debug_overlay.playerY\[-2\] _05107_ _05110_ rbzero.debug_overlay.playerY\[-3\]
+ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__a221o_1
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _09595_ _09596_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__nor2_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13718_ _06812_ _06813_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__xnor2_1
X_17486_ _01775_ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__and2b_1
X_14698_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__buf_4
XFILLER_176_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16437_ _08327_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__clkbuf_4
X_19225_ rbzero.spi_registers.new_texadd\[2\]\[9\] _03206_ _03220_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00840_ sky130_fd_sc_hd__o211a_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _06732_ _06727_ _06735_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__or3b_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19156_ rbzero.spi_registers.texadd1\[4\] _03176_ vssd1 vssd1 vccd1 vccd1 _03181_
+ sky130_fd_sc_hd__or2_1
X_16368_ _09457_ _09459_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ _09859_ _02385_ _02340_ rbzero.wall_tracer.trackDistY\[-4\] vssd1 vssd1 vccd1
+ vccd1 _00557_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_185_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15319_ _08390_ _08409_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__nor2_1
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19087_ rbzero.spi_registers.got_new_texadd\[0\] _03096_ vssd1 vssd1 vccd1 vccd1
+ _03140_ sky130_fd_sc_hd__nand2_2
X_16299_ _09146_ _08620_ _09389_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__o21ai_1
X_18038_ _02273_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20000_ _03639_ _03642_ _03584_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19989_ _03632_ _03633_ _03561_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21951_ net477 _01540_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ clknet_leaf_53_i_clk _00491_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21882_ net408 _01471_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20833_ clknet_leaf_67_i_clk _00422_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20764_ _09749_ _02747_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__and3_1
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20695_ _03908_ _03909_ _03910_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__nand3_1
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20291__157 clknet_1_0__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__inv_2
XFILLER_164_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21316_ clknet_leaf_31_i_clk _00905_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21247_ clknet_leaf_26_i_clk _00836_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ rbzero.tex_b1\[36\] rbzero.tex_b1\[37\] _04292_ vssd1 vssd1 vccd1 vccd1 _04298_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21178_ clknet_leaf_13_i_clk _00767_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20129_ _04589_ _05283_ _03721_ _04408_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a31o_1
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ rbzero.wall_tracer.mapX\[9\] rbzero.wall_tracer.mapX\[8\] rbzero.wall_tracer.mapX\[10\]
+ rbzero.wall_tracer.mapY\[7\] vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__or4_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ _05075_ _05080_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__o21ai_1
X_15670_ _08726_ _08753_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12882_ _06046_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__and2_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _07672_ _07791_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__xnor2_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _05021_ _05022_ _04819_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _10179_ _10233_ _10231_ vssd1 vssd1 vccd1 vccd1 _10359_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14552_ _07640_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__xor2_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _04947_ _04949_ _04951_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__o211a_1
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _06647_ _06673_ _06666_ _06598_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__a22o_1
XFILLER_201_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17271_ _08152_ _08399_ _10289_ vssd1 vssd1 vccd1 vccd1 _10290_ sky130_fd_sc_hd__or3_1
X_10715_ _04148_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14483_ _07417_ _07204_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__nor2_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ _04834_ _04884_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a21oi_1
X_19010_ _03090_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__clkbuf_1
X_16222_ _09053_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13434_ _06480_ _06482_ _06603_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__mux2_1
X_10646_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _04110_ vssd1 vssd1 vccd1 vccd1 _04112_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16153_ _09130_ _09132_ _09245_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__a21bo_1
XFILLER_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _06535_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__inv_2
X_10577_ _04075_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20350__210 clknet_1_0__leaf__03788_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__inv_2
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _08160_ _08198_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__nor2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ rbzero.tex_b0\[42\] _04913_ _04817_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a21o_1
X_16084_ _08410_ _08447_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__or2_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13296_ _06459_ _06461_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nor3_4
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19912_ rbzero.pov.ready_buffer\[64\] _03438_ _03558_ _03575_ vssd1 vssd1 vccd1 vccd1
+ _03576_ sky130_fd_sc_hd__a211o_1
X_15035_ rbzero.mapdyw\[1\] _06159_ _06255_ _08131_ vssd1 vssd1 vccd1 vccd1 _08132_
+ sky130_fd_sc_hd__a22o_1
X_12247_ rbzero.tex_g1\[57\] _04891_ _05031_ _04917_ vssd1 vssd1 vccd1 vccd1 _05434_
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19843_ _03533_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
X_12178_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _04932_ vssd1 vssd1 vccd1 vccd1 _05366_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11129_ _04365_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__clkbuf_1
X_19774_ _03497_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
X_16986_ _09587_ _09590_ _09719_ vssd1 vssd1 vccd1 vccd1 _10008_ sky130_fd_sc_hd__a21o_1
XFILLER_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18725_ _02914_ _02918_ _02915_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a21bo_1
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15937_ _09026_ _09031_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15868_ _08960_ _08962_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__xor2_1
X_18656_ rbzero.wall_tracer.rayAddendY\[4\] _02858_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02859_ sky130_fd_sc_hd__mux2_1
XFILLER_184_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17607_ rbzero.wall_tracer.visualWallDist\[5\] _08421_ vssd1 vssd1 vccd1 vccd1 _01898_
+ sky130_fd_sc_hd__nand2_1
X_14819_ _06595_ _07977_ _07978_ _07979_ _06631_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__a311o_1
X_15799_ _08887_ _08892_ _08893_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18587_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__clkbuf_4
X_17538_ _09542_ _09560_ _01722_ _01829_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__o31ai_1
XFILLER_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17469_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__nor2_1
XFILLER_149_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19208_ rbzero.spi_registers.texadd2\[2\] _03208_ vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19139_ rbzero.spi_registers.new_texadd\[0\]\[21\] _03140_ _03170_ _03169_ vssd1
+ vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__o211a_1
XFILLER_69_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21101_ clknet_leaf_72_i_clk _00690_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21032_ clknet_leaf_15_i_clk _00621_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_2
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19680__59 clknet_1_1__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21934_ net460 _01523_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21865_ net391 _01454_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ clknet_leaf_61_i_clk _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_21796_ net322 _01385_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20747_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
XFILLER_184_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ rbzero.tex_r1\[15\] rbzero.tex_r1\[16\] _04024_ vssd1 vssd1 vccd1 vccd1 _04033_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11480_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__clkinv_2
X_20678_ rbzero.texV\[5\] _03814_ _03819_ _03897_ vssd1 vssd1 vccd1 vccd1 _01616_
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10431_ rbzero.tex_r1\[48\] rbzero.tex_r1\[49\] _03991_ vssd1 vssd1 vccd1 vccd1 _03997_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__or2_1
XFILLER_136_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ _05279_ _05282_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21bo_1
XFILLER_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _06233_ _06248_ _06256_ _06142_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__a31o_2
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12032_ rbzero.tex_r1\[27\] _05195_ _05220_ _04923_ vssd1 vssd1 vccd1 vccd1 _05221_
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _09863_ _09864_ vssd1 vssd1 vccd1 vccd1 _09865_ sky130_fd_sc_hd__nor2_1
XFILLER_24_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16771_ _08942_ _08988_ _09803_ vssd1 vssd1 vccd1 vccd1 _09804_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13983_ _07108_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15722_ _08213_ _08297_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__or2_1
X_18510_ _09866_ _09767_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__or3_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12934_ _04679_ rbzero.map_rom.f4 _06107_ rbzero.debug_overlay.playerY\[3\] _06109_
+ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a221o_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19490_ rbzero.spi_registers.new_mapd\[9\] rbzero.spi_registers.spi_buffer\[9\] _03361_
+ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__mux2_1
XFILLER_160_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _08728_ _08747_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__xor2_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _02655_ _02656_ _02658_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__and3_1
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12865_ _06039_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or2_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _07773_ _07774_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__and2_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _04909_ vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__mux2_1
X_18372_ _02588_ _02604_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15584_ _08670_ _08678_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__and2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12796_ _05946_ _05968_ _05970_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a31o_1
XFILLER_57_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _10341_ vssd1 vssd1 vccd1 vccd1 _10342_ sky130_fd_sc_hd__clkbuf_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _07685_ _07705_ _07703_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__a21oi_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _04890_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__buf_6
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17254_ _10182_ _10199_ vssd1 vssd1 vccd1 vccd1 _10273_ sky130_fd_sc_hd__or2b_1
XFILLER_175_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__05700_ clknet_0__05700_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05700_
+ sky130_fd_sc_hd__clkbuf_16
X_14466_ _07630_ _07633_ _07635_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__nand3_1
X_11678_ rbzero.row_render.size\[6\] _04418_ _04867_ gpout0.hpos\[7\] vssd1 vssd1
+ vccd1 vccd1 _04868_ sky130_fd_sc_hd__o22a_1
XFILLER_179_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16205_ _09292_ _09181_ _09297_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__o21ai_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _06356_ _06481_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__xor2_1
X_10629_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _04099_ vssd1 vssd1 vccd1 vccd1 _04103_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17185_ _10080_ _10089_ vssd1 vssd1 vccd1 vccd1 _10205_ sky130_fd_sc_hd__and2b_1
XFILLER_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397_ _07558_ _07563_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__nand2_1
XFILLER_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16136_ _09103_ _09101_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__and2b_1
X_13348_ _06486_ _06492_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nand2_1
XFILLER_155_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ _09150_ _09160_ vssd1 vssd1 vccd1 vccd1 _09161_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _06393_ _06406_ _06411_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__a21oi_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15018_ _08119_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19826_ rbzero.pov.spi_buffer\[50\] rbzero.pov.spi_buffer\[51\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
XFILLER_111_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19757_ _03488_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
X_16969_ _09661_ _09704_ _09990_ vssd1 vssd1 vccd1 vccd1 _09991_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18708_ _02794_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__inv_2
X_19688_ clknet_1_0__leaf__03457_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__buf_1
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18639_ _02841_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__nand2_1
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21650_ clknet_leaf_85_i_clk _01239_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20322__186 clknet_1_1__leaf__03784_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__inv_2
XFILLER_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20601_ _03830_ _03831_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21581_ clknet_leaf_70_i_clk _01170_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22064_ clknet_leaf_79_i_clk _01653_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21015_ clknet_leaf_77_i_clk _00604_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10980_ _04287_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21917_ net443 _01506_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ net24 vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__buf_2
X_21848_ net374 _01437_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ _04772_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__nor2_1
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20297__163 clknet_1_1__leaf__03782_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__inv_2
X_12581_ reg_gpout\[1\] clknet_1_1__leaf__05761_ _05058_ vssd1 vssd1 vccd1 vccd1 _05762_
+ sky130_fd_sc_hd__mux2_2
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21779_ net305 _01368_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14320_ _07306_ _07208_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__nor2_1
XFILLER_184_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11532_ _04720_ _03973_ _04578_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a22o_1
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14251_ _07367_ _07368_ _07420_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__a21o_1
XFILLER_172_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ _04652_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13202_ _06370_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__or2_1
XFILLER_183_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10414_ rbzero.tex_r1\[56\] rbzero.tex_r1\[57\] _03980_ vssd1 vssd1 vccd1 vccd1 _03988_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14182_ _07347_ _07351_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__and2_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _04512_ _04477_ _04510_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__and3_1
XFILLER_48_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__nand2_1
X_18990_ _02474_ rbzero.spi_registers.spi_cmd\[0\] _03078_ vssd1 vssd1 vccd1 vccd1
+ _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_155_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17941_ _02137_ _02228_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__xnor2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ rbzero.map_overlay.i_otherx\[1\] _06117_ _06228_ rbzero.map_overlay.i_otherx\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a22o_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12015_ rbzero.tex_r1\[1\] _04982_ _05032_ _04919_ vssd1 vssd1 vccd1 vccd1 _05204_
+ sky130_fd_sc_hd__a31o_1
X_17872_ _02090_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__nand2_1
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20462__311 clknet_1_1__leaf__03799_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__inv_2
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19611_ _03434_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
X_16823_ _09839_ _09841_ _09840_ vssd1 vssd1 vccd1 vccd1 _09850_ sky130_fd_sc_hd__a21boi_1
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19542_ _03399_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__clkbuf_1
X_20557__17 clknet_1_0__leaf__03808_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
X_13966_ _07133_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__and2_1
XFILLER_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16754_ rbzero.wall_tracer.mapX\[8\] _09119_ vssd1 vssd1 vccd1 vccd1 _09790_ sky130_fd_sc_hd__xor2_1
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ _08796_ _08799_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__nand2_1
X_12917_ _06086_ _06076_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19473_ _03363_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
X_16685_ rbzero.row_render.size\[8\] _09752_ _09754_ _07992_ vssd1 vssd1 vccd1 vccd1
+ _00491_ sky130_fd_sc_hd__a22o_1
X_13897_ _07067_ _06741_ _07066_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__a21oi_1
XFILLER_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _02596_ _05106_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__or2_1
XFILLER_206_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15636_ _08233_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__clkbuf_4
X_12848_ _06019_ _06020_ _06022_ _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o211a_1
XFILLER_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ _08646_ _08647_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__xnor2_1
X_18355_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__and2_1
X_12779_ net40 _05944_ _05941_ net51 _05952_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a221o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ _10322_ _10324_ vssd1 vssd1 vccd1 vccd1 _10325_ sky130_fd_sc_hd__xor2_1
X_14518_ _07678_ _07688_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15498_ _08267_ _08288_ _08266_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__a21bo_1
X_18286_ rbzero.wall_tracer.rayAddendX\[-5\] _02523_ _02525_ vssd1 vssd1 vccd1 vccd1
+ _02526_ sky130_fd_sc_hd__mux2_1
XFILLER_147_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17237_ _10255_ _10256_ vssd1 vssd1 vccd1 vccd1 _10257_ sky130_fd_sc_hd__nand2_1
X_14449_ _07602_ _07618_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__nor2_1
XFILLER_163_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ _10186_ _10187_ vssd1 vssd1 vccd1 vccd1 _10188_ sky130_fd_sc_hd__and2_1
XFILLER_157_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16119_ _09024_ _09067_ _09212_ vssd1 vssd1 vccd1 vccd1 _09213_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17099_ _10118_ _10119_ vssd1 vssd1 vccd1 vccd1 _10120_ sky130_fd_sc_hd__nor2_2
XFILLER_157_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19809_ rbzero.pov.spi_buffer\[42\] rbzero.pov.spi_buffer\[43\] _03512_ vssd1 vssd1
+ vccd1 vccd1 _03516_ sky130_fd_sc_hd__mux2_1
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21702_ net228 _01291_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21633_ clknet_leaf_79_i_clk _01222_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21564_ clknet_leaf_92_i_clk _01153_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21495_ net213 _01084_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20446_ clknet_1_1__leaf__03796_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__buf_1
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22047_ clknet_leaf_55_i_clk _01636_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _06990_ _06943_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ _06914_ _06915_ _06921_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__nor3_1
XFILLER_44_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10963_ _04278_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12702_ _05880_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20305__170 clknet_1_0__leaf__03783_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__inv_2
X_16470_ _08950_ _09560_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__nor2_1
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13682_ _06785_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__nor2_1
XFILLER_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _04242_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _08265_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12633_ _05797_ _05800_ _05805_ _05812_ _05793_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a32o_2
XFILLER_106_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ _08149_ _08445_ _08446_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__a21oi_2
X_18140_ _02411_ _02412_ _02413_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__and3_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ _05055_ _05719_ _05720_ net71 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a22o_1
XFILLER_200_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14303_ _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__or2_1
XFILLER_157_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18071_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__nand2_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ rbzero.map_overlay.i_otherx\[2\] vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__inv_2
X_15283_ _06073_ _06349_ rbzero.side_hot vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__mux2_1
X_12495_ _05642_ _05657_ _05676_ net8 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__o22ai_1
X_17022_ _09519_ _08618_ _09079_ _09520_ vssd1 vssd1 vccd1 vccd1 _10043_ sky130_fd_sc_hd__o22ai_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14234_ _07341_ _07355_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__nor2_1
X_11446_ _04445_ _04448_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__nor2_4
XFILLER_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _07264_ _07290_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__or2b_1
XFILLER_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ _04454_ _04534_ _04540_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or3_1
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] _06286_
+ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nand3_1
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18973_ rbzero.spi_registers.spi_buffer\[17\] rbzero.spi_registers.spi_buffer\[16\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _06640_ _06769_ _06720_ _06722_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__o22a_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _02210_ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__nor2_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _06088_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__nand2_1
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _02136_ _02047_ _02142_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__and3_1
XFILLER_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _09825_ _09827_ _09826_ vssd1 vssd1 vccd1 vccd1 _09835_ sky130_fd_sc_hd__a21boi_1
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17786_ _01878_ _02075_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14998_ rbzero.wall_tracer.stepDistX\[4\] _08012_ _08103_ vssd1 vssd1 vccd1 vccd1
+ _08109_ sky130_fd_sc_hd__mux2_1
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19525_ _03390_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
X_16737_ _06129_ _09118_ vssd1 vssd1 vccd1 vccd1 _09775_ sky130_fd_sc_hd__xnor2_1
X_13949_ _06741_ _07066_ _07069_ _07070_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__a22o_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19456_ rbzero.spi_registers.new_vshift\[2\] _02483_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03354_ sky130_fd_sc_hd__mux2_1
X_16668_ _04051_ _04637_ _05053_ _09727_ vssd1 vssd1 vccd1 vccd1 _09747_ sky130_fd_sc_hd__and4_1
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18407_ _02635_ _02636_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nand2_1
X_15619_ _08227_ _08276_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__nor2_1
XFILLER_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19387_ _03314_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16599_ _08148_ _09688_ _08454_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__a21o_1
X_18338_ _02568_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18269_ _02509_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21280_ clknet_leaf_1_i_clk _00869_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469__317 clknet_1_0__leaf__03800_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__inv_2
XFILLER_162_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03789_ clknet_0__03789_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03789_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20162_ _05652_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__inv_2
XFILLER_104_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20093_ rbzero.pov.ready_buffer\[20\] _03684_ _03700_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01228_ sky130_fd_sc_hd__o211a_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20995_ clknet_leaf_0_i_clk _00584_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21616_ clknet_leaf_90_i_clk _01205_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21547_ clknet_leaf_92_i_clk _01136_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ rbzero.spi_registers.texadd0\[7\] _04466_ _04490_ _04491_ vssd1 vssd1 vccd1
+ vccd1 _04492_ sky130_fd_sc_hd__o22a_1
XFILLER_193_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _04702_ _05462_ _05464_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a31oi_1
XFILLER_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21478_ net196 _01067_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ _04426_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_4
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11162_ _04382_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15970_ _08480_ _08493_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__or2b_1
X_11093_ _04346_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14921_ _04442_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__buf_2
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _01929_ _01930_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__xor2_1
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14852_ _06577_ _07826_ _07871_ _06631_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__a31o_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _06790_ _06687_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__nor2_1
X_17571_ _01766_ _01750_ _01861_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14783_ _06641_ _07902_ _06670_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11995_ rbzero.tex_r1\[15\] _04933_ _05183_ _04923_ vssd1 vssd1 vccd1 vccd1 _05184_
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19310_ rbzero.spi_registers.texadd3\[22\] _03241_ vssd1 vssd1 vccd1 vccd1 _03269_
+ sky130_fd_sc_hd__or2_1
X_16522_ _09539_ _09518_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__or2b_1
XFILLER_21_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13734_ _06761_ _06904_ _06748_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10946_ _04269_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19241_ rbzero.spi_registers.texadd2\[16\] _03222_ vssd1 vssd1 vccd1 vccd1 _03230_
+ sky130_fd_sc_hd__or2_1
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16453_ _09293_ _09410_ _09543_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__a21bo_1
X_13665_ _06742_ _06743_ _06640_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__a21o_1
X_10877_ _04233_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _08424_ _08427_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__and2_2
X_12616_ net19 _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
XFILLER_169_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19172_ rbzero.spi_registers.new_texadd\[1\]\[10\] _03188_ _03190_ _03184_ vssd1
+ vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__o211a_1
X_16384_ _09121_ _09474_ _09475_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__a21o_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _06378_ _06544_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__nand2_2
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15335_ _08410_ _08390_ _08400_ _08429_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__or4_1
X_18123_ _09873_ _02399_ _02340_ rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1
+ vccd1 _00559_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _05724_ _05725_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__o21a_1
XFILLER_184_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _08346_ _08356_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_144_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18054_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__buf_2
XFILLER_144_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ _05055_ _05637_ _05659_ net71 vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a22oi_1
XANTENNA_3 _04464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _09910_ _09924_ _10025_ vssd1 vssd1 vccd1 vccd1 _10026_ sky130_fd_sc_hd__a21o_1
X_14217_ _07385_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11429_ rbzero.spi_registers.texadd1\[2\] _04545_ _04536_ _04620_ vssd1 vssd1 vccd1
+ vccd1 _04621_ sky130_fd_sc_hd__a211o_1
X_15197_ rbzero.wall_tracer.stepDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__inv_2
XFILLER_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14148_ _07305_ _07315_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__o21a_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18956_ rbzero.spi_registers.spi_buffer\[9\] rbzero.spi_registers.spi_buffer\[8\]
+ _03052_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
X_14079_ _06720_ _07249_ _07204_ _07206_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__o22ai_1
XFILLER_112_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _01718_ _02194_ _02106_ _02107_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a2bb2o_1
X_18887_ rbzero.pov.spi_buffer\[51\] rbzero.pov.ready_buffer\[51\] _03022_ vssd1 vssd1
+ vccd1 vccd1 _03025_ sky130_fd_sc_hd__mux2_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17838_ _02125_ _02126_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nand2_1
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17769_ _02043_ _02058_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__xor2_1
X_20223__96 clknet_1_1__leaf__03465_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19508_ rbzero.spi_registers.got_new_texadd\[0\] _08117_ _03316_ _03381_ vssd1 vssd1
+ vccd1 vccd1 _00962_ sky130_fd_sc_hd__a31o_1
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20780_ gpout2.clk_div\[0\] net63 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_1
X_20440__291 clknet_1_1__leaf__03797_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__inv_2
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _03344_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21401_ clknet_leaf_28_i_clk _00990_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21332_ clknet_leaf_31_i_clk _00921_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21263_ clknet_leaf_3_i_clk _00852_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20214_ rbzero.spi_registers.new_texadd\[3\]\[22\] rbzero.spi_registers.spi_buffer\[22\]
+ _03384_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux2_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21194_ clknet_leaf_29_i_clk _00783_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20145_ _09732_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__buf_4
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03801_ clknet_0__03801_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03801_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ rbzero.pov.ready_buffer\[12\] _03684_ _03691_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01220_ sky130_fd_sc_hd__o211a_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ rbzero.tex_g1\[3\] rbzero.tex_g1\[4\] _04188_ vssd1 vssd1 vccd1 vccd1 _04193_
+ sky130_fd_sc_hd__mux2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _04914_ vssd1 vssd1 vccd1 vccd1 _04970_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20978_ clknet_leaf_63_i_clk _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ rbzero.tex_g1\[36\] rbzero.tex_g1\[37\] _04155_ vssd1 vssd1 vccd1 vccd1 _04157_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _06486_ _06492_ _06603_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__mux2_1
X_10662_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _04110_ vssd1 vssd1 vccd1 vccd1 _04120_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _05190_ _05583_ _05585_ _04952_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__o211a_1
XFILLER_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ _06463_ _06551_ _06448_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__o21a_1
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10593_ rbzero.tex_r0\[38\] rbzero.tex_r0\[37\] _04077_ vssd1 vssd1 vccd1 vccd1 _04084_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ rbzero.debug_overlay.playerX\[-6\] _08207_ vssd1 vssd1 vccd1 vccd1 _08215_
+ sky130_fd_sc_hd__or2_1
X_20417__271 clknet_1_1__leaf__03794_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__inv_2
X_12332_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _04908_ vssd1 vssd1 vccd1 vccd1 _05518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19686__65 clknet_1_0__leaf__03461_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
X_15051_ _04430_ _08141_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__or2_1
XFILLER_108_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ rbzero.tex_g1\[34\] _04830_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or2_1
XFILLER_135_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14002_ _07169_ _07172_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__inv_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12194_ _04429_ _04635_ _05056_ _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__o211a_4
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__buf_2
X_18810_ _02984_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
Xoutput73 net125 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__clkbuf_1
X_11145_ rbzero.tex_b0\[32\] rbzero.tex_b0\[31\] _04373_ vssd1 vssd1 vccd1 vccd1 _04374_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19790_ rbzero.pov.spi_buffer\[33\] rbzero.pov.spi_buffer\[34\] _03501_ vssd1 vssd1
+ vccd1 vccd1 _03506_ sky130_fd_sc_hd__mux2_1
XFILLER_62_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18741_ _02475_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o21ai_1
XFILLER_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11076_ _04337_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
X_15953_ _08462_ _08465_ _08458_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__a21oi_2
XFILLER_23_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14904_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.trackDistX\[-8\] _08037_
+ vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__mux2_1
X_18672_ _02854_ _02872_ _02867_ _04434_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a31o_1
XFILLER_209_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _08973_ _08974_ _08976_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__o21bai_1
XFILLER_23_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _01893_ _01913_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__xnor2_2
XFILLER_64_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14835_ _06575_ _07813_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__nand2_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _01843_ _01844_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__and2_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ rbzero.debug_overlay.playerY\[4\] _05095_ _05096_ rbzero.debug_overlay.playerY\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__a22o_1
X_14766_ _07928_ _07930_ _07932_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__a21o_1
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16505_ _09593_ _09594_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__and2_1
X_10929_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _04259_ vssd1 vssd1 vccd1 vccd1 _04261_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13717_ _06782_ _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__xnor2_1
X_17485_ _09519_ _09242_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or3_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _04436_ _04437_ _04433_ _06259_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__and4b_2
XFILLER_205_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19224_ rbzero.spi_registers.texadd2\[9\] _03208_ vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__or2_1
X_16436_ _09524_ _09526_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13648_ _06765_ _06817_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__nor3b_1
XFILLER_13_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19155_ rbzero.spi_registers.new_texadd\[1\]\[3\] _03174_ _03180_ _03169_ vssd1 vssd1
+ vccd1 vccd1 _00810_ sky130_fd_sc_hd__o211a_1
X_16367_ _09267_ _09332_ _09458_ vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13579_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__nor2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18106_ _02383_ _02384_ _02337_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__o21a_1
X_15318_ _08410_ _08400_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__nor2_1
X_16298_ _09146_ _08553_ _09389_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__or3_1
XFILLER_184_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19086_ rbzero.spi_registers.new_mapd\[1\] _03119_ _03139_ _03130_ vssd1 vssd1 vccd1
+ vccd1 _00782_ sky130_fd_sc_hd__o211a_1
XFILLER_184_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037_ _02321_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _08343_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_68_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ rbzero.debug_overlay.playerY\[0\] _08320_ vssd1 vssd1 vccd1 vccd1 _03633_
+ sky130_fd_sc_hd__nand2_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18939_ _03053_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21950_ net476 _01539_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
X_20245__116 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__inv_2
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20901_ clknet_leaf_53_i_clk _00490_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21881_ net407 _01470_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20832_ clknet_leaf_67_i_clk _00421_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_165_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20763_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__or2_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20694_ _03908_ _03909_ _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__a21o_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21315_ clknet_leaf_31_i_clk _00904_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21246_ clknet_leaf_26_i_clk _00835_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21177_ clknet_leaf_20_i_clk _00766_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20128_ _04698_ _04413_ _03977_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__and3b_1
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20447__297 clknet_1_1__leaf__03798_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__inv_2
X_12950_ rbzero.wall_tracer.mapX\[5\] vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__inv_2
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ rbzero.pov.ready_buffer\[27\] _03656_ _03680_ _03681_ vssd1 vssd1 vccd1 vccd1
+ _01213_ sky130_fd_sc_hd__o211a_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _05080_ _05082_ _05085_ _05086_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a41o_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _06010_ _06017_ _06005_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a21o_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\] vssd1 vssd1 vccd1
+ vccd1 _05022_ sky130_fd_sc_hd__nand2_1
X_14620_ _07671_ _07713_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nor2_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14551_ _07252_ _07476_ _07721_ _07719_ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__o31a_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11763_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__buf_6
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ rbzero.tex_g1\[44\] rbzero.tex_g1\[45\] _04144_ vssd1 vssd1 vccd1 vccd1 _04148_
+ sky130_fd_sc_hd__mux2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _06512_ _06603_ _06586_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__a21o_1
XFILLER_187_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17270_ _10288_ _08428_ vssd1 vssd1 vccd1 vccd1 _10289_ sky130_fd_sc_hd__or2_1
X_14482_ _07611_ _07610_ _07609_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__a21o_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11694_ rbzero.row_render.size\[10\] rbzero.row_render.size\[9\] _04841_ _04883_
+ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__or4_2
XFILLER_201_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16221_ _08466_ _09184_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__nand2_1
X_13433_ _06455_ _06461_ _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__mux2_1
X_10645_ _04111_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _09008_ _08618_ _09077_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__or3_1
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13364_ _06530_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nand2_1
X_10576_ rbzero.tex_r0\[46\] rbzero.tex_r0\[45\] _04066_ vssd1 vssd1 vccd1 vccd1 _04075_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ rbzero.tex_b0\[43\] _04926_ _04928_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__and3_1
XFILLER_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15103_ _04463_ _06056_ _08143_ _08197_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__o211a_1
X_16083_ _08434_ _09176_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__nor2_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13295_ _06463_ _06465_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__or2_1
X_19911_ _08256_ _03570_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__nor2_1
X_15034_ _06159_ _08126_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__nor2_1
X_12246_ rbzero.tex_g1\[59\] _04964_ _05432_ _04946_ vssd1 vssd1 vccd1 vccd1 _05433_
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19842_ rbzero.pov.spi_buffer\[58\] rbzero.pov.spi_buffer\[59\] _03523_ vssd1 vssd1
+ vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
X_12177_ rbzero.tex_g0\[63\] _04927_ _04929_ _05199_ vssd1 vssd1 vccd1 vccd1 _05365_
+ sky130_fd_sc_hd__a31o_1
XFILLER_64_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11128_ rbzero.tex_b0\[40\] rbzero.tex_b0\[39\] _04362_ vssd1 vssd1 vccd1 vccd1 _04365_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19773_ rbzero.pov.spi_buffer\[25\] rbzero.pov.spi_buffer\[26\] _03490_ vssd1 vssd1
+ vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
X_16985_ _09720_ vssd1 vssd1 vccd1 vccd1 _10007_ sky130_fd_sc_hd__inv_2
XFILLER_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18724_ rbzero.wall_tracer.rayAddendY\[9\] _02525_ _09760_ _02919_ _02921_ vssd1
+ vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__o221a_1
XFILLER_83_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15936_ _09029_ _09030_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__xor2_1
X_11059_ rbzero.tex_b1\[8\] rbzero.tex_b1\[9\] _04325_ vssd1 vssd1 vccd1 vccd1 _04329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18655_ _08134_ _02852_ _02856_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__o22a_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _08344_ _08950_ _08954_ _08961_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__o31a_1
XFILLER_97_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17606_ _10315_ _09252_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__or2_1
XFILLER_149_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14818_ _06595_ _07950_ vssd1 vssd1 vccd1 vccd1 _07979_ sky130_fd_sc_hd__nor2_1
XFILLER_149_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _09753_ _02789_ _02790_ _02793_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__a31o_1
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15798_ _08871_ _08886_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__and2b_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17537_ _08889_ _01718_ _01720_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__or3_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14749_ _07827_ _07872_ _07871_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__a21o_1
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17468_ _06170_ _09785_ _01760_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19207_ rbzero.spi_registers.new_texadd\[2\]\[1\] _03206_ _03210_ _03197_ vssd1 vssd1
+ vccd1 vccd1 _00832_ sky130_fd_sc_hd__o211a_1
X_16419_ _09495_ _09509_ vssd1 vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__xnor2_1
X_17399_ _10386_ _01691_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19138_ rbzero.spi_registers.texadd0\[21\] _03142_ vssd1 vssd1 vccd1 vccd1 _03170_
+ sky130_fd_sc_hd__or2_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19069_ rbzero.map_overlay.i_mapdy\[1\] _03122_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__or2_1
XFILLER_106_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21100_ clknet_leaf_71_i_clk _00689_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19665__46 clknet_1_1__leaf__03459_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21031_ clknet_leaf_46_i_clk _00620_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_2
XFILLER_114_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21933_ net459 _01522_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21864_ net390 _01453_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20815_ clknet_leaf_61_i_clk _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21795_ net321 _01384_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20746_ gpout0.clk_div\[0\] net63 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nor2_1
XFILLER_168_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20677_ _03893_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10430_ _03996_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _04653_ _04695_ _05284_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__o2111a_1
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__inv_2
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ rbzero.tex_r1\[26\] _05032_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__or2_1
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21229_ clknet_leaf_2_i_clk _00818_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20529__372 clknet_1_1__leaf__03805_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__inv_2
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20228__100 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__inv_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16770_ _08942_ _08988_ _08123_ vssd1 vssd1 vccd1 vccd1 _09803_ sky130_fd_sc_hd__a21oi_1
X_13982_ _07148_ _07152_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__xnor2_1
X_20380__237 clknet_1_1__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__inv_2
XFILLER_111_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15721_ _08516_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__clkbuf_4
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ rbzero.debug_overlay.playerX\[0\] _06108_ rbzero.map_rom.i_row\[4\] _04673_
+ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a22o_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _02656_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__inv_2
X_15652_ _08743_ _08746_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__and2_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _05996_ _05998_ _06029_ _06038_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__and4_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _07771_ _07772_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__nand2_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _04920_ _04999_ _05004_ _04902_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a211o_1
X_18371_ _02602_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15583_ _08670_ _08676_ _08677_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__nand3_1
X_12795_ _05946_ _05971_ net37 vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17322_ _10340_ _10092_ _10331_ vssd1 vssd1 vccd1 vccd1 _10341_ sky130_fd_sc_hd__or3b_1
XFILLER_144_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ rbzero.tex_r0\[2\] _04933_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a21o_1
X_14534_ _07703_ _07704_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nor2_1
XFILLER_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17253_ _10159_ _10176_ _10174_ vssd1 vssd1 vccd1 vccd1 _10272_ sky130_fd_sc_hd__a21o_1
XFILLER_144_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14465_ _07630_ _07633_ _07635_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__a21o_1
X_11677_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] vssd1 vssd1 vccd1
+ vccd1 _04867_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20274__142 clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__inv_2
X_16204_ _09295_ _09296_ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__xnor2_1
X_10628_ _04102_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13416_ _06545_ _06558_ _06564_ _06474_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__o31a_1
X_17184_ _09974_ _09975_ _08910_ vssd1 vssd1 vccd1 vccd1 _10204_ sky130_fd_sc_hd__a21o_1
X_14396_ _07565_ _07566_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13347_ _06408_ _06464_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__xor2_1
X_16135_ _09227_ _09228_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__xnor2_1
X_10559_ _04054_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ _09158_ _09159_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__nor2_1
X_13278_ _04444_ _06341_ _06343_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ rbzero.tex_g1\[25\] _04904_ _05182_ _04918_ vssd1 vssd1 vccd1 vccd1 _05416_
+ sky130_fd_sc_hd__a31o_1
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15017_ _08117_ _05382_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__and2_1
XFILLER_68_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19825_ _03524_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19756_ rbzero.pov.spi_buffer\[17\] rbzero.pov.spi_buffer\[18\] _03479_ vssd1 vssd1
+ vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
X_16968_ _09701_ _09703_ vssd1 vssd1 vccd1 vccd1 _09990_ sky130_fd_sc_hd__and2b_1
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18707_ _02903_ _02904_ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21oi_1
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15919_ _09012_ _09013_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16899_ _09911_ _09920_ vssd1 vssd1 vccd1 vccd1 _09921_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18638_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nand2_1
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18569_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__nand2_1
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20600_ _03825_ _03828_ _03826_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a21boi_1
XFILLER_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21580_ clknet_leaf_70_i_clk _01169_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_opt_4_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22063_ clknet_leaf_79_i_clk _01652_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21014_ clknet_leaf_77_i_clk _00603_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21916_ net442 _01505_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21847_ net373 _01436_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11600_ _04778_ _04786_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__o21a_1
XFILLER_12_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12580_ _05710_ _05759_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__a21oi_2
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21778_ net304 _01367_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ rbzero.map_overlay.i_mapdx\[1\] vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__inv_2
X_20729_ _03728_ clknet_1_0__leaf__05938_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__and2_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14250_ _07367_ _07368_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__nand3_1
X_11462_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__buf_4
XFILLER_165_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13201_ rbzero.wall_tracer.rayAddendX\[-2\] _06371_ _06323_ vssd1 vssd1 vccd1 vccd1
+ _06372_ sky130_fd_sc_hd__mux2_2
XFILLER_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10413_ _03987_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__clkbuf_1
X_14181_ _07347_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nor2_1
XFILLER_165_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11393_ _04518_ _04520_ _04462_ _04517_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a211oi_1
XFILLER_109_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ _06299_ _06300_ _06301_ _06302_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__o211a_1
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17940_ _02007_ _09315_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__nor2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _06237_ _06144_ _06130_ rbzero.map_overlay.i_othery\[0\] _06238_ vssd1 vssd1
+ vccd1 vccd1 _06239_ sky130_fd_sc_hd__a221o_1
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12014_ rbzero.tex_r1\[3\] _05195_ _05202_ _04923_ vssd1 vssd1 vccd1 vccd1 _05203_
+ sky130_fd_sc_hd__o211a_1
X_17871_ _02158_ _02159_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__xor2_1
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19610_ rbzero.spi_registers.new_texadd\[1\]\[22\] rbzero.spi_registers.spi_buffer\[22\]
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16822_ _09847_ _09848_ vssd1 vssd1 vccd1 vccd1 _09849_ sky130_fd_sc_hd__or2b_1
XFILLER_171_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19541_ rbzero.spi_registers.new_texadd\[0\]\[12\] rbzero.spi_registers.spi_buffer\[12\]
+ _03395_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
X_16753_ rbzero.wall_tracer.mapX\[7\] _09786_ _09784_ _09789_ vssd1 vssd1 vccd1 vccd1
+ _00524_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13965_ _06687_ _06769_ _07135_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _08796_ _08797_ _08798_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__nand3_1
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12916_ rbzero.map_rom.c6 _06077_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a21o_1
X_19472_ rbzero.spi_registers.new_mapd\[0\] _02473_ _03362_ vssd1 vssd1 vccd1 vccd1
+ _03363_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16684_ _09753_ vssd1 vssd1 vccd1 vccd1 _09754_ sky130_fd_sc_hd__buf_4
X_13896_ _06767_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__buf_4
X_18423_ _02635_ _02641_ _02650_ _08134_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a31o_1
XFILLER_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ _08201_ _08440_ _08665_ _08667_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12847_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nand2_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__nor2_1
XFILLER_15_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15566_ _08652_ _08660_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__nand2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ net46 _05944_ _05953_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a211o_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _09397_ _09037_ _10191_ _10323_ vssd1 vssd1 vccd1 vccd1 _10324_ sky130_fd_sc_hd__o31a_1
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _07252_ _07444_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nor2_1
X_11729_ _04918_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__clkbuf_8
X_18285_ _02524_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__buf_4
X_15497_ _08513_ _08574_ _08591_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__a21o_1
XFILLER_175_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _10009_ _10249_ _10252_ vssd1 vssd1 vccd1 vccd1 _10256_ sky130_fd_sc_hd__o21a_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14448_ _07602_ _07618_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__xor2_1
XFILLER_190_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17167_ _10059_ _08620_ _10185_ vssd1 vssd1 vccd1 vccd1 _10187_ sky130_fd_sc_hd__o21ai_1
XFILLER_155_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14379_ _07362_ _07445_ _07479_ _07549_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__o211a_1
XFILLER_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16118_ _09064_ _09066_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__nor2_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10119_ sky130_fd_sc_hd__and2_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16049_ _09083_ _09142_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19808_ _03515_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19739_ _03467_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21701_ net227 _01290_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21632_ clknet_leaf_80_i_clk _01221_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21563_ clknet_leaf_92_i_clk _01152_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21494_ net212 _01083_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20411__266 clknet_1_1__leaf__03793_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__inv_2
XFILLER_133_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22046_ clknet_leaf_55_i_clk _01635_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ rbzero.tex_b1\[54\] rbzero.tex_b1\[55\] _04270_ vssd1 vssd1 vccd1 vccd1 _04278_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13750_ _06919_ _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__nand2_1
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12701_ reg_gpout\[3\] clknet_1_0__leaf__05879_ net45 vssd1 vssd1 vccd1 vccd1 _05880_
+ sky130_fd_sc_hd__mux2_2
XFILLER_189_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10893_ rbzero.tex_g0\[24\] rbzero.tex_g0\[23\] _04237_ vssd1 vssd1 vccd1 vccd1 _04242_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13681_ _06830_ _06831_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nor2_1
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15420_ _08496_ _08514_ vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__xor2_1
X_12632_ _05765_ _05770_ _05807_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a31o_2
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20492__338 clknet_1_0__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__inv_2
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15351_ rbzero.wall_tracer.stepDistX\[2\] _08357_ _08405_ rbzero.wall_tracer.stepDistY\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__a22o_1
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _05707_ _05739_ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__or3_1
XFILLER_15_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11514_ _04411_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__buf_4
X_14302_ _07464_ _07462_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__xor2_2
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18070_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__or2_1
X_15282_ _08368_ _08265_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__nor2_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ _05660_ _05662_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__o21ba_1
XFILLER_138_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17021_ _09936_ _09938_ vssd1 vssd1 vccd1 vccd1 _10042_ sky130_fd_sc_hd__nand2_1
X_14233_ _07402_ _07403_ _07396_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__a21oi_1
X_11445_ net2 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__clkinv_2
XFILLER_109_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _07333_ _07334_ _06540_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11376_ _04452_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or2_1
XFILLER_4_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13115_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__or2_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18972_ _03070_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__clkbuf_1
X_14095_ _07264_ _07265_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__nand2_1
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20386__243 clknet_1_0__leaf__03791_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__inv_2
X_17923_ _02186_ _02116_ _02209_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__nor3_1
XFILLER_117_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _06144_ _06088_ _06218_ _06221_ rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1
+ _06222_ sky130_fd_sc_hd__a221o_1
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17854_ _02136_ _02047_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16805_ _09832_ _09833_ vssd1 vssd1 vccd1 vccd1 _09834_ sky130_fd_sc_hd__or2b_1
XFILLER_208_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17785_ _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nor2_1
XFILLER_208_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14997_ _08108_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19524_ rbzero.spi_registers.new_texadd\[0\]\[4\] _02487_ _03381_ vssd1 vssd1 vccd1
+ vccd1 _03390_ sky130_fd_sc_hd__mux2_1
X_16736_ _09765_ _09772_ _09773_ vssd1 vssd1 vccd1 vccd1 _09774_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13948_ _07117_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__and2_1
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19455_ _03353_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16667_ _09745_ vssd1 vssd1 vccd1 vccd1 _09746_ sky130_fd_sc_hd__buf_4
X_13879_ _07036_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__and2b_1
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18406_ _02596_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02636_
+ sky130_fd_sc_hd__or2_1
X_15618_ _08672_ _08712_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__xor2_1
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19386_ _02487_ rbzero.spi_registers.new_sky\[4\] _03309_ vssd1 vssd1 vccd1 vccd1
+ _03314_ sky130_fd_sc_hd__mux2_1
X_16598_ _08027_ _08029_ _08031_ _09563_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__or4_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18337_ _02570_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__or2_1
X_15549_ _08635_ _08640_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__nor2_1
XFILLER_33_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18268_ rbzero.spi_registers.new_texadd\[2\]\[23\] rbzero.spi_registers.spi_buffer\[23\]
+ _02478_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _10146_ _10238_ vssd1 vssd1 vccd1 vccd1 _10239_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18199_ _02456_ _02458_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03788_ clknet_0__03788_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03788_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20161_ _03745_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20092_ _02681_ _03655_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ clknet_leaf_1_i_clk _00583_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21615_ clknet_leaf_90_i_clk _01204_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21546_ clknet_leaf_90_i_clk _01135_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_127_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21477_ net195 _01066_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _03975_ _04417_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a21boi_2
XFILLER_181_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19701__78 clknet_1_0__leaf__03463_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ rbzero.tex_b0\[24\] rbzero.tex_b0\[23\] _04373_ vssd1 vssd1 vccd1 vccd1 _04382_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _04340_ vssd1 vssd1 vccd1 vccd1 _04346_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22029_ clknet_leaf_55_i_clk _01618_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_1
X_14920_ rbzero.wall_tracer.visualWallDist\[-3\] _08047_ vssd1 vssd1 vccd1 vccd1 _08060_
+ sky130_fd_sc_hd__or2_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ _08007_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13802_ _06969_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__and2b_1
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17570_ _01766_ _01750_ _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__and3_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14782_ _07894_ _07926_ _07946_ _06641_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__o211a_1
X_11994_ rbzero.tex_r1\[14\] _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or2_1
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16521_ _09495_ _09509_ _09507_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__a21o_1
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13733_ _06658_ _06725_ _06756_ _06760_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a22o_1
X_10945_ rbzero.tex_b1\[62\] rbzero.tex_b1\[63\] _04188_ vssd1 vssd1 vccd1 vccd1 _04269_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19240_ rbzero.spi_registers.new_texadd\[2\]\[15\] _03221_ _03229_ _03226_ vssd1
+ vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__o211a_1
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16452_ _09542_ _08497_ _09411_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__or3_1
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13664_ _06750_ _06733_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__nor2_1
X_10876_ rbzero.tex_g0\[32\] rbzero.tex_g0\[31\] _04226_ vssd1 vssd1 vccd1 vccd1 _04233_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15403_ _08497_ _08441_ _08487_ _08488_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__a2bb2o_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ net49 _05791_ _05792_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__o2bb2a_1
X_19171_ rbzero.spi_registers.texadd1\[10\] _03189_ vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__or2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _09121_ _09474_ _08145_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__o21ai_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _06740_ _06752_ _06753_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__a31o_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _02341_ _02397_ _02398_ _02337_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__o31a_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _08420_ _06263_ _08421_ _08422_ _08428_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__o221a_2
X_12546_ _05711_ _05726_ _05712_ net15 vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a31o_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18053_ _02336_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__buf_4
X_15265_ _08328_ _08337_ _08343_ _08325_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__o22a_1
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ net5 _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nor2_1
XFILLER_184_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17004_ _09921_ _09923_ vssd1 vssd1 vccd1 vccd1 _10025_ sky130_fd_sc_hd__nor2_1
XFILLER_172_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_4 _04464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _07347_ _07386_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__and2_1
X_11428_ rbzero.spi_registers.texadd2\[2\] _04537_ _04457_ rbzero.spi_registers.texadd3\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a22o_1
X_15196_ _08246_ _08253_ _08265_ _08276_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__o22ai_1
XFILLER_153_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11359_ rbzero.spi_registers.texadd1\[21\] _04545_ _04536_ _04550_ vssd1 vssd1 vccd1
+ vccd1 _04551_ sky130_fd_sc_hd__a211o_1
X_14147_ _07316_ _07249_ _07317_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__or3b_1
XFILLER_28_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14078_ _07248_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__clkbuf_4
X_18955_ _03061_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17906_ _08530_ _02105_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__nand2_1
X_13029_ rbzero.wall_tracer.trackDistX\[1\] _06199_ _06204_ vssd1 vssd1 vccd1 vccd1
+ _06205_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18886_ _03024_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17837_ _10315_ _09363_ _02124_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17768_ _02049_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16719_ rbzero.traced_texa\[10\] _09759_ _09758_ rbzero.wall_tracer.visualWallDist\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a22o_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19507_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__buf_4
X_17699_ _01986_ _01987_ _09866_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a21o_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19438_ rbzero.spi_registers.spi_buffer\[6\] rbzero.spi_registers.new_other\[6\]
+ _03338_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__mux2_1
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19369_ rbzero.spi_registers.vshift\[4\] _03298_ vssd1 vssd1 vccd1 vccd1 _03304_
+ sky130_fd_sc_hd__or2_1
XFILLER_163_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21400_ clknet_leaf_6_i_clk _00989_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21331_ clknet_leaf_31_i_clk _00920_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21262_ clknet_leaf_3_i_clk _00851_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20213_ _03773_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21193_ clknet_leaf_22_i_clk _00782_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20144_ _03716_ _03729_ _03733_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a21oi_1
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03800_ clknet_0__03800_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03800_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20075_ rbzero.debug_overlay.vplaneX\[-8\] _03685_ vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__or2_1
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20977_ clknet_leaf_63_i_clk _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10730_ _04156_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _04119_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12400_ _05198_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
XFILLER_185_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13380_ _06499_ _06489_ _06523_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__o31ai_1
X_10592_ _04083_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _05515_ _05516_ _04934_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__mux2_1
XFILLER_182_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21529_ clknet_leaf_97_i_clk _01118_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12262_ rbzero.tex_g1\[36\] _04904_ _04964_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_
+ sky130_fd_sc_hd__a31o_1
X_15050_ _08144_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__clkbuf_8
XFILLER_177_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11213_ _04409_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_8
X_14001_ _07170_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__and2b_1
XFILLER_108_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12193_ _05051_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__nand2_1
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ _04214_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__clkbuf_4
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 o_reset sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__buf_2
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18740_ rbzero.spi_registers.spi_cmd\[0\] _02474_ vssd1 vssd1 vccd1 vccd1 _02936_
+ sky130_fd_sc_hd__and2_1
XFILLER_62_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15952_ _09044_ _09046_ _08441_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__a21oi_2
X_11075_ rbzero.tex_b1\[0\] rbzero.tex_b1\[1\] _03979_ vssd1 vssd1 vccd1 vccd1 _04337_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14903_ _08036_ _08044_ _08048_ _01633_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__o211a_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18671_ _02854_ _02867_ _02872_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a21oi_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08935_ _08977_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__and2_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _01911_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__nor2_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _07993_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20498__344 clknet_1_0__leaf__03802_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__inv_2
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ _01843_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__nor2_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _06669_ _07931_ _06470_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__a21o_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11977_ rbzero.debug_overlay.playerY\[-9\] _05122_ _05118_ rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a22o_1
XFILLER_189_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16504_ _09593_ _09594_ vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__nor2_1
XFILLER_205_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13716_ _06850_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10928_ _04260_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
X_17484_ _09647_ _09362_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__or2_1
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14696_ _06470_ _07865_ _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__o21ai_4
XFILLER_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19223_ rbzero.spi_registers.new_texadd\[2\]\[8\] _03206_ _03219_ _03213_ vssd1 vssd1
+ vccd1 vccd1 _00839_ sky130_fd_sc_hd__o211a_1
XFILLER_189_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16435_ _09525_ _08620_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13647_ _06803_ _06815_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__xor2_1
X_10859_ rbzero.tex_g0\[40\] rbzero.tex_g0\[39\] _04215_ vssd1 vssd1 vccd1 vccd1 _04224_
+ sky130_fd_sc_hd__mux2_1
XFILLER_176_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ rbzero.spi_registers.texadd1\[3\] _03176_ vssd1 vssd1 vccd1 vccd1 _03180_
+ sky130_fd_sc_hd__or2_1
X_16366_ _09329_ _09331_ vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__nor2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13578_ _06682_ _06693_ _06700_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ _02380_ _02381_ _02382_ _06104_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a31o_1
X_15317_ _08228_ _08384_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__or2_1
XFILLER_121_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19085_ rbzero.mapdyw\[1\] _03121_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__or2_1
X_12529_ _05702_ _05703_ net15 _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__or4_1
X_16297_ _09387_ _09388_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__nand2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18036_ _02243_ _02244_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__o21a_1
X_15248_ rbzero.wall_tracer.stepDistX\[-10\] _06263_ _08159_ _08163_ vssd1 vssd1 vccd1
+ vccd1 _08343_ sky130_fd_sc_hd__o22ai_4
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ rbzero.wall_tracer.stepDistY\[-7\] _08157_ _08270_ _08273_ vssd1 vssd1 vccd1
+ vccd1 _08274_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19987_ rbzero.debug_overlay.playerY\[0\] _08320_ vssd1 vssd1 vccd1 vccd1 _03632_
+ sky130_fd_sc_hd__or2_1
XFILLER_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18938_ _02473_ rbzero.spi_registers.mosi _03052_ vssd1 vssd1 vccd1 vccd1 _03053_
+ sky130_fd_sc_hd__mux2_1
.ends


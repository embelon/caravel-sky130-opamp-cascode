// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net73;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net74;
 wire net89;
 wire net90;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net107;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.otherx[0] ;
 wire \rbzero.otherx[1] ;
 wire \rbzero.otherx[2] ;
 wire \rbzero.otherx[3] ;
 wire \rbzero.otherx[4] ;
 wire \rbzero.othery[0] ;
 wire \rbzero.othery[1] ;
 wire \rbzero.othery[2] ;
 wire \rbzero.othery[3] ;
 wire \rbzero.othery[4] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.texu[5] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-12] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[11] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[11] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-12] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[11] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[11] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[11] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[11] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[11] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.side ;
 wire \rbzero.wall_tracer.state[0] ;
 wire \rbzero.wall_tracer.state[10] ;
 wire \rbzero.wall_tracer.state[11] ;
 wire \rbzero.wall_tracer.state[12] ;
 wire \rbzero.wall_tracer.state[13] ;
 wire \rbzero.wall_tracer.state[14] ;
 wire \rbzero.wall_tracer.state[1] ;
 wire \rbzero.wall_tracer.state[2] ;
 wire \rbzero.wall_tracer.state[3] ;
 wire \rbzero.wall_tracer.state[4] ;
 wire \rbzero.wall_tracer.state[5] ;
 wire \rbzero.wall_tracer.state[6] ;
 wire \rbzero.wall_tracer.state[7] ;
 wire \rbzero.wall_tracer.state[8] ;
 wire \rbzero.wall_tracer.state[9] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-12] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[11] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-12] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[11] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.texu[0] ;
 wire \rbzero.wall_tracer.texu[1] ;
 wire \rbzero.wall_tracer.texu[2] ;
 wire \rbzero.wall_tracer.texu[3] ;
 wire \rbzero.wall_tracer.texu[4] ;
 wire \rbzero.wall_tracer.texu[5] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-12] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[11] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-12] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[11] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-12] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[11] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \rbzero.wall_tracer.wall[0] ;
 wire \rbzero.wall_tracer.wall[1] ;
 wire net91;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_leaf_0_i_clk;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net126;
 wire net71;
 wire net72;
 wire net123;
 wire net124;
 wire net125;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_2_0_i_clk;
 wire clknet_opt_3_0_i_clk;
 wire clknet_opt_4_0_i_clk;
 wire clknet_opt_5_0_i_clk;
 wire clknet_opt_6_0_i_clk;
 wire clknet_opt_6_1_i_clk;
 wire clknet_opt_7_0_i_clk;
 wire clknet_opt_8_0_i_clk;
 wire clknet_opt_9_0_i_clk;
 wire clknet_opt_10_0_i_clk;
 wire clknet_opt_10_1_i_clk;
 wire clknet_opt_11_0_i_clk;
 wire clknet_opt_12_0_i_clk;
 wire clknet_opt_13_0_i_clk;
 wire clknet_0__04835_;
 wire clknet_1_0__leaf__04835_;
 wire clknet_1_1__leaf__04835_;
 wire clknet_0__03321_;
 wire clknet_1_0__leaf__03321_;
 wire clknet_1_1__leaf__03321_;
 wire clknet_0__03320_;
 wire clknet_1_0__leaf__03320_;
 wire clknet_1_1__leaf__03320_;
 wire clknet_0__03309_;
 wire clknet_1_0__leaf__03309_;
 wire clknet_1_1__leaf__03309_;
 wire clknet_0__03319_;
 wire clknet_1_0__leaf__03319_;
 wire clknet_1_1__leaf__03319_;
 wire clknet_0__03318_;
 wire clknet_1_0__leaf__03318_;
 wire clknet_1_1__leaf__03318_;
 wire clknet_0__03317_;
 wire clknet_1_0__leaf__03317_;
 wire clknet_1_1__leaf__03317_;
 wire clknet_0__03316_;
 wire clknet_1_0__leaf__03316_;
 wire clknet_1_1__leaf__03316_;
 wire clknet_0__03315_;
 wire clknet_1_0__leaf__03315_;
 wire clknet_1_1__leaf__03315_;
 wire clknet_0__03314_;
 wire clknet_1_0__leaf__03314_;
 wire clknet_1_1__leaf__03314_;
 wire clknet_0__03313_;
 wire clknet_1_0__leaf__03313_;
 wire clknet_1_1__leaf__03313_;
 wire clknet_0__03312_;
 wire clknet_1_0__leaf__03312_;
 wire clknet_1_1__leaf__03312_;
 wire clknet_0__03311_;
 wire clknet_1_0__leaf__03311_;
 wire clknet_1_1__leaf__03311_;
 wire clknet_0__03310_;
 wire clknet_1_0__leaf__03310_;
 wire clknet_1_1__leaf__03310_;
 wire clknet_0__03298_;
 wire clknet_1_0__leaf__03298_;
 wire clknet_1_1__leaf__03298_;
 wire clknet_0__03308_;
 wire clknet_1_0__leaf__03308_;
 wire clknet_1_1__leaf__03308_;
 wire clknet_0__03307_;
 wire clknet_1_0__leaf__03307_;
 wire clknet_1_1__leaf__03307_;
 wire clknet_0__03306_;
 wire clknet_1_0__leaf__03306_;
 wire clknet_1_1__leaf__03306_;
 wire clknet_0__03305_;
 wire clknet_1_0__leaf__03305_;
 wire clknet_1_1__leaf__03305_;
 wire clknet_0__03304_;
 wire clknet_1_0__leaf__03304_;
 wire clknet_1_1__leaf__03304_;
 wire clknet_0__03303_;
 wire clknet_1_0__leaf__03303_;
 wire clknet_1_1__leaf__03303_;
 wire clknet_0__03302_;
 wire clknet_1_0__leaf__03302_;
 wire clknet_1_1__leaf__03302_;
 wire clknet_0__03301_;
 wire clknet_1_0__leaf__03301_;
 wire clknet_1_1__leaf__03301_;
 wire clknet_0__03300_;
 wire clknet_1_0__leaf__03300_;
 wire clknet_1_1__leaf__03300_;
 wire clknet_0__03299_;
 wire clknet_1_0__leaf__03299_;
 wire clknet_1_1__leaf__03299_;
 wire clknet_0__03044_;
 wire clknet_1_0__leaf__03044_;
 wire clknet_1_1__leaf__03044_;
 wire clknet_0__03297_;
 wire clknet_1_0__leaf__03297_;
 wire clknet_1_1__leaf__03297_;
 wire clknet_0__03296_;
 wire clknet_1_0__leaf__03296_;
 wire clknet_1_1__leaf__03296_;
 wire clknet_0__03295_;
 wire clknet_1_0__leaf__03295_;
 wire clknet_1_1__leaf__03295_;
 wire clknet_0__03294_;
 wire clknet_1_0__leaf__03294_;
 wire clknet_1_1__leaf__03294_;
 wire clknet_0__03293_;
 wire clknet_1_0__leaf__03293_;
 wire clknet_1_1__leaf__03293_;
 wire clknet_0__03292_;
 wire clknet_1_0__leaf__03292_;
 wire clknet_1_1__leaf__03292_;
 wire clknet_0__03291_;
 wire clknet_1_0__leaf__03291_;
 wire clknet_1_1__leaf__03291_;
 wire clknet_0__03290_;
 wire clknet_1_0__leaf__03290_;
 wire clknet_1_1__leaf__03290_;
 wire clknet_0__03289_;
 wire clknet_1_0__leaf__03289_;
 wire clknet_1_1__leaf__03289_;
 wire clknet_0__03045_;
 wire clknet_1_0__leaf__03045_;
 wire clknet_1_1__leaf__03045_;
 wire clknet_0__03037_;
 wire clknet_1_0__leaf__03037_;
 wire clknet_1_1__leaf__03037_;
 wire clknet_0__03043_;
 wire clknet_1_0__leaf__03043_;
 wire clknet_1_1__leaf__03043_;
 wire clknet_0__03042_;
 wire clknet_1_0__leaf__03042_;
 wire clknet_1_1__leaf__03042_;
 wire clknet_0__03041_;
 wire clknet_1_0__leaf__03041_;
 wire clknet_1_1__leaf__03041_;
 wire clknet_0__03040_;
 wire clknet_1_0__leaf__03040_;
 wire clknet_1_1__leaf__03040_;
 wire clknet_0__03039_;
 wire clknet_1_0__leaf__03039_;
 wire clknet_1_1__leaf__03039_;
 wire clknet_0__03038_;
 wire clknet_1_0__leaf__03038_;
 wire clknet_1_1__leaf__03038_;
 wire net54;
 wire net70;
 wire net511;
 wire net512;
 wire net513;
 wire net514;

 sky130_fd_sc_hd__buf_4 _10298_ (.A(\gpout0.hpos[0] ),
    .X(_03473_));
 sky130_fd_sc_hd__buf_4 _10299_ (.A(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__buf_4 _10300_ (.A(\gpout0.hpos[7] ),
    .X(_03475_));
 sky130_fd_sc_hd__inv_2 _10301_ (.A(\gpout0.hpos[8] ),
    .Y(_03476_));
 sky130_fd_sc_hd__clkbuf_4 _10302_ (.A(\gpout0.hpos[9] ),
    .X(_03477_));
 sky130_fd_sc_hd__and2_1 _10303_ (.A(_03476_),
    .B(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__xor2_4 _10304_ (.A(net45),
    .B(net44),
    .X(_03479_));
 sky130_fd_sc_hd__buf_6 _10305_ (.A(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__and4_1 _10306_ (.A(_03474_),
    .B(_03475_),
    .C(_03478_),
    .D(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_4 _10307_ (.A(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_4 _10308_ (.A(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net46),
    .S(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _10310_ (.A(_03484_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10311_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_03483_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_1 _10312_ (.A(_03485_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _10313_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_03483_),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_1 _10314_ (.A(_03486_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_03483_),
    .X(_03487_));
 sky130_fd_sc_hd__clkbuf_1 _10316_ (.A(_03487_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10317_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_03483_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _10318_ (.A(_03488_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_03483_),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_1 _10320_ (.A(_03489_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_03483_),
    .X(_03490_));
 sky130_fd_sc_hd__clkbuf_1 _10322_ (.A(_03490_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10323_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_03483_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_1 _10324_ (.A(_03491_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _10325_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_03483_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _10326_ (.A(_03492_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10327_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_03483_),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_1 _10328_ (.A(_03493_),
    .X(_01372_));
 sky130_fd_sc_hd__clkbuf_4 _10329_ (.A(_03482_),
    .X(_03494_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_1 _10331_ (.A(_03495_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10332_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_03494_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_1 _10333_ (.A(_03496_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_03494_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_1 _10335_ (.A(_03497_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_03494_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_1 _10337_ (.A(_03498_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10338_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_03494_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _10339_ (.A(_03499_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10340_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_03494_),
    .X(_03500_));
 sky130_fd_sc_hd__clkbuf_1 _10341_ (.A(_03500_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_03494_),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_1 _10343_ (.A(_03501_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_03494_),
    .X(_03502_));
 sky130_fd_sc_hd__clkbuf_1 _10345_ (.A(_03502_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_03494_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_1 _10347_ (.A(_03503_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10348_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_03494_),
    .X(_03504_));
 sky130_fd_sc_hd__clkbuf_1 _10349_ (.A(_03504_),
    .X(_01362_));
 sky130_fd_sc_hd__clkbuf_4 _10350_ (.A(_03482_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _10351_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _10352_ (.A(_03506_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_03505_),
    .X(_03507_));
 sky130_fd_sc_hd__clkbuf_1 _10354_ (.A(_03507_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _10355_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_03505_),
    .X(_03508_));
 sky130_fd_sc_hd__clkbuf_1 _10356_ (.A(_03508_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _10357_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_03505_),
    .X(_03509_));
 sky130_fd_sc_hd__clkbuf_1 _10358_ (.A(_03509_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(\rbzero.tex_r1[39] ),
    .A1(net54),
    .S(_03505_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_1 _10360_ (.A(_03510_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_03505_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _10362_ (.A(_03511_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10363_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_03505_),
    .X(_03512_));
 sky130_fd_sc_hd__clkbuf_1 _10364_ (.A(_03512_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10365_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_03505_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_1 _10366_ (.A(_03513_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_03505_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_1 _10368_ (.A(_03514_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_03505_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _10370_ (.A(_03515_),
    .X(_01352_));
 sky130_fd_sc_hd__clkbuf_4 _10371_ (.A(_03482_),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_1 _10372_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__clkbuf_1 _10373_ (.A(_03517_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10374_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_03516_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _10375_ (.A(_03518_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _10376_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_03516_),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_1 _10377_ (.A(_03519_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10378_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_03516_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_1 _10379_ (.A(_03520_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10380_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_03516_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_1 _10381_ (.A(_03521_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10382_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_03516_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _10383_ (.A(_03522_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10384_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_03516_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _10385_ (.A(_03523_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10386_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_03516_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _10387_ (.A(_03524_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_03516_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _10389_ (.A(_03525_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10390_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_03516_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _10391_ (.A(_03526_),
    .X(_01342_));
 sky130_fd_sc_hd__clkbuf_4 _10392_ (.A(_03482_),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_1 _10393_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _10394_ (.A(_03528_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10395_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_03527_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _10396_ (.A(_03529_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _10397_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_03527_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _10398_ (.A(_03530_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _10399_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_03527_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _10400_ (.A(_03531_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _10401_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_03527_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _10402_ (.A(_03532_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _10403_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_03527_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _10404_ (.A(_03533_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _10405_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_03527_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _10406_ (.A(_03534_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _10407_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_03527_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _10408_ (.A(_03535_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _10409_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_03527_),
    .X(_03536_));
 sky130_fd_sc_hd__clkbuf_1 _10410_ (.A(_03536_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _10411_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_03527_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _10412_ (.A(_03537_),
    .X(_01332_));
 sky130_fd_sc_hd__clkbuf_4 _10413_ (.A(_03482_),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_03539_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_03538_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_03540_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_03538_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _10419_ (.A(_03541_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_03538_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _10421_ (.A(_03542_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_03538_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _10423_ (.A(_03543_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_03538_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _10425_ (.A(_03544_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_03538_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _10427_ (.A(_03545_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_03538_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _10429_ (.A(_03546_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _10430_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_03538_),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _10431_ (.A(_03547_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_03538_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _10433_ (.A(_03548_),
    .X(_01322_));
 sky130_fd_sc_hd__clkbuf_4 _10434_ (.A(_03482_),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _10436_ (.A(_03550_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_03551_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_03549_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _10440_ (.A(_03552_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_03549_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _10442_ (.A(_03553_),
    .X(_01318_));
 sky130_fd_sc_hd__nand2_2 _10443_ (.A(_03475_),
    .B(_03478_),
    .Y(_03554_));
 sky130_fd_sc_hd__inv_12 _10444_ (.A(_03479_),
    .Y(_03555_));
 sky130_fd_sc_hd__or3_2 _10445_ (.A(_03474_),
    .B(_03554_),
    .C(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_4 _10446_ (.A(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__clkbuf_4 _10447_ (.A(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(net46),
    .A1(\rbzero.tex_r0[63] ),
    .S(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _10449_ (.A(_03559_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _10450_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_03558_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _10451_ (.A(_03560_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _10452_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_03558_),
    .X(_03561_));
 sky130_fd_sc_hd__clkbuf_1 _10453_ (.A(_03561_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_03558_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _10455_ (.A(_03562_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_03558_),
    .X(_03563_));
 sky130_fd_sc_hd__clkbuf_1 _10457_ (.A(_03563_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_03558_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _10459_ (.A(_03564_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_03558_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_03565_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_03558_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _10463_ (.A(_03566_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_03558_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _10465_ (.A(_03567_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_03558_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_1 _10467_ (.A(_03568_),
    .X(_01308_));
 sky130_fd_sc_hd__clkbuf_4 _10468_ (.A(_03557_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(_03570_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_03569_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _10472_ (.A(_03571_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_03569_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _10474_ (.A(_03572_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_03569_),
    .X(_03573_));
 sky130_fd_sc_hd__clkbuf_1 _10476_ (.A(_03573_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_03569_),
    .X(_03574_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_03574_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_03569_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_1 _10480_ (.A(_03575_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_03569_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_03576_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_03569_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_1 _10484_ (.A(_03577_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_03569_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_03578_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_03569_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_03579_),
    .X(_01298_));
 sky130_fd_sc_hd__clkbuf_4 _10489_ (.A(_03557_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_1 _10491_ (.A(_03581_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_03580_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _10493_ (.A(_03582_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_03580_),
    .X(_03583_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_03583_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_03580_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _10497_ (.A(_03584_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_03580_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_03585_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_03580_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _10501_ (.A(_03586_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _10502_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_03580_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _10503_ (.A(_03587_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_03580_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _10505_ (.A(_03588_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_03580_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _10507_ (.A(_03589_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_03580_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _10509_ (.A(_03590_),
    .X(_01288_));
 sky130_fd_sc_hd__clkbuf_4 _10510_ (.A(_03557_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _10512_ (.A(_03592_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_03591_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _10514_ (.A(_03593_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_03591_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _10516_ (.A(_03594_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_03591_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _10518_ (.A(_03595_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_03591_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _10520_ (.A(_03596_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_03591_),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _10522_ (.A(_03597_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _10523_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_03591_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _10524_ (.A(_03598_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_03591_),
    .X(_03599_));
 sky130_fd_sc_hd__clkbuf_1 _10526_ (.A(_03599_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_03591_),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _10528_ (.A(_03600_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_03591_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _10530_ (.A(_03601_),
    .X(_01278_));
 sky130_fd_sc_hd__clkbuf_4 _10531_ (.A(_03557_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _10533_ (.A(_03603_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_03602_),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_1 _10535_ (.A(_03604_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_03602_),
    .X(_03605_));
 sky130_fd_sc_hd__clkbuf_1 _10537_ (.A(_03605_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_03602_),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_1 _10539_ (.A(_03606_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_03602_),
    .X(_03607_));
 sky130_fd_sc_hd__clkbuf_1 _10541_ (.A(_03607_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_03602_),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _10543_ (.A(_03608_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _10544_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_03602_),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_1 _10545_ (.A(_03609_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_03602_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_03610_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_03602_),
    .X(_03611_));
 sky130_fd_sc_hd__clkbuf_1 _10549_ (.A(_03611_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_03602_),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _10551_ (.A(_03612_),
    .X(_01268_));
 sky130_fd_sc_hd__clkbuf_4 _10552_ (.A(_03557_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_1 _10554_ (.A(_03614_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_03613_),
    .X(_03615_));
 sky130_fd_sc_hd__clkbuf_1 _10556_ (.A(_03615_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_03613_),
    .X(_03616_));
 sky130_fd_sc_hd__clkbuf_1 _10558_ (.A(_03616_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_03613_),
    .X(_03617_));
 sky130_fd_sc_hd__clkbuf_1 _10560_ (.A(_03617_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_03613_),
    .X(_03618_));
 sky130_fd_sc_hd__clkbuf_1 _10562_ (.A(_03618_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_03613_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _10564_ (.A(_03619_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _10565_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_03613_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _10566_ (.A(_03620_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_03613_),
    .X(_03621_));
 sky130_fd_sc_hd__clkbuf_1 _10568_ (.A(_03621_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_03613_),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_1 _10570_ (.A(_03622_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_03613_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_03623_),
    .X(_01258_));
 sky130_fd_sc_hd__clkbuf_4 _10573_ (.A(_03557_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_1 _10575_ (.A(_03625_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_03624_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _10577_ (.A(_03626_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_03624_),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_1 _10579_ (.A(_03627_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_03624_),
    .X(_03628_));
 sky130_fd_sc_hd__clkbuf_1 _10581_ (.A(_03628_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net47),
    .S(_03549_),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _10583_ (.A(_03629_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _10584_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_03549_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_1 _10585_ (.A(_03630_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_03549_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _10587_ (.A(_03631_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_03549_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _10589_ (.A(_03632_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_03549_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_03633_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_03549_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_1 _10593_ (.A(_03634_),
    .X(_01248_));
 sky130_fd_sc_hd__clkbuf_4 _10594_ (.A(_03482_),
    .X(_03635_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_1 _10596_ (.A(_03636_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_03635_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _10598_ (.A(_03637_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_03635_),
    .X(_03638_));
 sky130_fd_sc_hd__clkbuf_1 _10600_ (.A(_03638_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_03635_),
    .X(_03639_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_03639_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_03635_),
    .X(_03640_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_03640_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_03635_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_03641_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_03635_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_03642_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_03635_),
    .X(_03643_));
 sky130_fd_sc_hd__clkbuf_1 _10610_ (.A(_03643_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_03635_),
    .X(_03644_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_03644_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_03635_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_03645_),
    .X(_01238_));
 sky130_fd_sc_hd__buf_4 _10615_ (.A(_03481_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_4 _10616_ (.A(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_1 _10618_ (.A(_03648_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_03647_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _10620_ (.A(_03649_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_03647_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_1 _10622_ (.A(_03650_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _10623_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_03647_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _10624_ (.A(_03651_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_03647_),
    .X(_03652_));
 sky130_fd_sc_hd__clkbuf_1 _10626_ (.A(_03652_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_03647_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_1 _10628_ (.A(_03653_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _10629_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_03647_),
    .X(_03654_));
 sky130_fd_sc_hd__clkbuf_1 _10630_ (.A(_03654_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_03647_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(_03655_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_03647_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _10634_ (.A(_03656_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_03647_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _10636_ (.A(_03657_),
    .X(_01228_));
 sky130_fd_sc_hd__clkbuf_4 _10637_ (.A(_03646_),
    .X(_03658_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_03659_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_03658_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_1 _10641_ (.A(_03660_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _10642_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_03658_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_1 _10643_ (.A(_03661_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_03658_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_1 _10645_ (.A(_03662_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_03658_),
    .X(_03663_));
 sky130_fd_sc_hd__clkbuf_1 _10647_ (.A(_03663_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_03658_),
    .X(_03664_));
 sky130_fd_sc_hd__clkbuf_1 _10649_ (.A(_03664_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_03658_),
    .X(_03665_));
 sky130_fd_sc_hd__clkbuf_1 _10651_ (.A(_03665_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_03658_),
    .X(_03666_));
 sky130_fd_sc_hd__clkbuf_1 _10653_ (.A(_03666_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_03658_),
    .X(_03667_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(_03667_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_03658_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _10657_ (.A(_03668_),
    .X(_01218_));
 sky130_fd_sc_hd__clkbuf_4 _10658_ (.A(_03646_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__clkbuf_1 _10660_ (.A(_03670_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_03669_),
    .X(_03671_));
 sky130_fd_sc_hd__clkbuf_1 _10662_ (.A(_03671_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_03669_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _10664_ (.A(_03672_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_03669_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _10666_ (.A(_03673_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _10667_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_03669_),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_1 _10668_ (.A(_03674_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_03669_),
    .X(_03675_));
 sky130_fd_sc_hd__clkbuf_1 _10670_ (.A(_03675_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _10671_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_03669_),
    .X(_03676_));
 sky130_fd_sc_hd__clkbuf_1 _10672_ (.A(_03676_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_03669_),
    .X(_03677_));
 sky130_fd_sc_hd__clkbuf_1 _10674_ (.A(_03677_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_03669_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _10676_ (.A(_03678_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _10677_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_03669_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_1 _10678_ (.A(_03679_),
    .X(_01208_));
 sky130_fd_sc_hd__clkbuf_4 _10679_ (.A(_03646_),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_03681_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_03680_),
    .X(_03682_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_03682_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_03680_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _10685_ (.A(_03683_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _10686_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_03680_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_1 _10687_ (.A(_03684_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_03680_),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_03685_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_03680_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _10691_ (.A(_03686_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_03680_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_1 _10693_ (.A(_03687_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_03680_),
    .X(_03688_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(_03688_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_03680_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(_03689_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_03680_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(_03690_),
    .X(_01198_));
 sky130_fd_sc_hd__clkbuf_4 _10700_ (.A(_03646_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_03692_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_03691_),
    .X(_03693_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_03693_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_03691_),
    .X(_03694_));
 sky130_fd_sc_hd__clkbuf_1 _10706_ (.A(_03694_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _10707_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_03691_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _10708_ (.A(_03695_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_03691_),
    .X(_03696_));
 sky130_fd_sc_hd__clkbuf_1 _10710_ (.A(_03696_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_03691_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_1 _10712_ (.A(_03697_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _10713_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_03691_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _10714_ (.A(_03698_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_03691_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_1 _10716_ (.A(_03699_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(net47),
    .A1(\rbzero.tex_g0[63] ),
    .S(_03624_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_1 _10718_ (.A(_03700_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_03624_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_1 _10720_ (.A(_03701_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_03624_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_1 _10722_ (.A(_03702_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_03624_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_1 _10724_ (.A(_03703_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_03624_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_03704_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_03624_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(_03705_),
    .X(_01184_));
 sky130_fd_sc_hd__clkbuf_4 _10729_ (.A(_03557_),
    .X(_03706_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_1 _10731_ (.A(_03707_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_03706_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_1 _10733_ (.A(_03708_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_03706_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_03709_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_03706_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(_03710_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_03706_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(_03711_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_03706_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(_03712_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_03706_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _10743_ (.A(_03713_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_03706_),
    .X(_03714_));
 sky130_fd_sc_hd__clkbuf_1 _10745_ (.A(_03714_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_03706_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(_03715_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_03706_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(_03716_),
    .X(_01174_));
 sky130_fd_sc_hd__buf_4 _10750_ (.A(_03556_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_4 _10751_ (.A(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(_03719_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_03718_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(_03720_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_03718_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(_03721_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_03718_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_03722_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_03718_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_03723_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_03718_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_03724_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_03718_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_03725_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_03718_),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_03726_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_03718_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_03727_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_03718_),
    .X(_03728_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(_03728_),
    .X(_01164_));
 sky130_fd_sc_hd__clkbuf_4 _10772_ (.A(_03717_),
    .X(_03729_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(_03730_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_03729_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(_03731_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_03729_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_03732_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_03729_),
    .X(_03733_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_03733_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_03729_),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_03734_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_03729_),
    .X(_03735_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_03735_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_03729_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_03736_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_03729_),
    .X(_03737_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(_03737_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_03729_),
    .X(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_03738_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_03729_),
    .X(_03739_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_03739_),
    .X(_01154_));
 sky130_fd_sc_hd__clkbuf_4 _10793_ (.A(_03717_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__clkbuf_1 _10795_ (.A(_03741_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_03740_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _10797_ (.A(_03742_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_03740_),
    .X(_03743_));
 sky130_fd_sc_hd__clkbuf_1 _10799_ (.A(_03743_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_03740_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(_03744_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_03740_),
    .X(_03745_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(_03745_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_03740_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(_03746_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_03740_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(_03747_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_03740_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(_03748_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_03740_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_03749_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_03740_),
    .X(_03750_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_03750_),
    .X(_01144_));
 sky130_fd_sc_hd__clkbuf_4 _10814_ (.A(_03717_),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _10816_ (.A(_03752_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_03751_),
    .X(_03753_));
 sky130_fd_sc_hd__clkbuf_1 _10818_ (.A(_03753_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_03751_),
    .X(_03754_));
 sky130_fd_sc_hd__clkbuf_1 _10820_ (.A(_03754_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_03751_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_03755_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_03751_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_03756_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_03751_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_03757_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_03751_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(_03758_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_03751_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_03759_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_03751_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_03760_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_03751_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_03761_),
    .X(_01134_));
 sky130_fd_sc_hd__buf_4 _10835_ (.A(_03717_),
    .X(_03762_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_1 _10837_ (.A(_03763_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_03762_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _10839_ (.A(_03764_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_03762_),
    .X(_03765_));
 sky130_fd_sc_hd__clkbuf_1 _10841_ (.A(_03765_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_03762_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _10843_ (.A(_03766_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_03762_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_1 _10845_ (.A(_03767_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_03762_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(_03768_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_03762_),
    .X(_03769_));
 sky130_fd_sc_hd__clkbuf_1 _10849_ (.A(_03769_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _10850_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_03762_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _10851_ (.A(_03770_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net48),
    .S(_03691_),
    .X(_03771_));
 sky130_fd_sc_hd__clkbuf_1 _10853_ (.A(_03771_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_03691_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _10855_ (.A(_03772_),
    .X(_01124_));
 sky130_fd_sc_hd__clkbuf_4 _10856_ (.A(_03646_),
    .X(_03773_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_03774_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_03773_),
    .X(_03775_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_03775_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_03773_),
    .X(_03776_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_03776_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_03773_),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(_03777_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_03773_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_1 _10866_ (.A(_03778_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_03773_),
    .X(_03779_));
 sky130_fd_sc_hd__clkbuf_1 _10868_ (.A(_03779_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_03773_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_1 _10870_ (.A(_03780_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_03773_),
    .X(_03781_));
 sky130_fd_sc_hd__clkbuf_1 _10872_ (.A(_03781_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_03773_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_1 _10874_ (.A(_03782_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_03773_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_1 _10876_ (.A(_03783_),
    .X(_01114_));
 sky130_fd_sc_hd__clkbuf_4 _10877_ (.A(_03646_),
    .X(_03784_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_03785_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_03784_),
    .X(_03786_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_03786_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_03784_),
    .X(_03787_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(_03787_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_03784_),
    .X(_03788_));
 sky130_fd_sc_hd__clkbuf_1 _10885_ (.A(_03788_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_03784_),
    .X(_03789_));
 sky130_fd_sc_hd__clkbuf_1 _10887_ (.A(_03789_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_03784_),
    .X(_03790_));
 sky130_fd_sc_hd__clkbuf_1 _10889_ (.A(_03790_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_03784_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_1 _10891_ (.A(_03791_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _10892_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_03784_),
    .X(_03792_));
 sky130_fd_sc_hd__clkbuf_1 _10893_ (.A(_03792_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _10894_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_03784_),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_1 _10895_ (.A(_03793_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _10896_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_03784_),
    .X(_03794_));
 sky130_fd_sc_hd__clkbuf_1 _10897_ (.A(_03794_),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_4 _10898_ (.A(_03646_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_03796_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_03795_),
    .X(_03797_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_03797_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_03795_),
    .X(_03798_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_03798_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_03795_),
    .X(_03799_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_03799_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_03795_),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_03800_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_03795_),
    .X(_03801_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_03801_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_03795_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_03802_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_03795_),
    .X(_03803_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_03803_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_03795_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_1 _10916_ (.A(_03804_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _10917_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_03795_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _10918_ (.A(_03805_),
    .X(_01094_));
 sky130_fd_sc_hd__clkbuf_4 _10919_ (.A(_03646_),
    .X(_03806_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(_03807_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_03806_),
    .X(_03808_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_03808_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_03806_),
    .X(_03809_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_03809_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_03806_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_03810_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_03806_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_03811_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_03806_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(_03812_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_03806_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _10933_ (.A(_03813_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _10934_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_03806_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _10935_ (.A(_03814_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_03806_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _10937_ (.A(_03815_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_03806_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _10939_ (.A(_03816_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_4 _10940_ (.A(_03646_),
    .X(_03817_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(_03818_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_03817_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_03819_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_03817_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_03820_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_03817_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_03821_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_03817_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_03822_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_03817_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(_03823_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_03817_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _10954_ (.A(_03824_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_03817_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_1 _10956_ (.A(_03825_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_03817_),
    .X(_03826_));
 sky130_fd_sc_hd__clkbuf_1 _10958_ (.A(_03826_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_03817_),
    .X(_03827_));
 sky130_fd_sc_hd__clkbuf_1 _10960_ (.A(_03827_),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_4 _10961_ (.A(_03481_),
    .X(_03828_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(_03829_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_03828_),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(_03830_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_03828_),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(_03831_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_03828_),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_03832_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_03828_),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_03833_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_03828_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_03834_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_03828_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(_03835_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_03828_),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _10977_ (.A(_03836_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_03828_),
    .X(_03837_));
 sky130_fd_sc_hd__clkbuf_1 _10979_ (.A(_03837_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_03828_),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_1 _10981_ (.A(_03838_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_03482_),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(_03839_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_03482_),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_03840_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(net48),
    .A1(\rbzero.tex_b0[63] ),
    .S(_03762_),
    .X(_03841_));
 sky130_fd_sc_hd__clkbuf_1 _10987_ (.A(_03841_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_03762_),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_1 _10989_ (.A(_03842_),
    .X(_00891_));
 sky130_fd_sc_hd__clkbuf_4 _10990_ (.A(_03717_),
    .X(_03843_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(_03844_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_03843_),
    .X(_03845_));
 sky130_fd_sc_hd__clkbuf_1 _10994_ (.A(_03845_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_03843_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _10996_ (.A(_03846_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_03843_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_1 _10998_ (.A(_03847_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_03843_),
    .X(_03848_));
 sky130_fd_sc_hd__clkbuf_1 _11000_ (.A(_03848_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_03843_),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_1 _11002_ (.A(_03849_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_03843_),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_03850_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_03843_),
    .X(_03851_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_03851_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_03843_),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(_03852_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_03843_),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(_03853_),
    .X(_00881_));
 sky130_fd_sc_hd__clkbuf_4 _11011_ (.A(_03717_),
    .X(_03854_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_1 _11013_ (.A(_03855_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_03854_),
    .X(_03856_));
 sky130_fd_sc_hd__clkbuf_1 _11015_ (.A(_03856_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_03854_),
    .X(_03857_));
 sky130_fd_sc_hd__clkbuf_1 _11017_ (.A(_03857_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_03854_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_1 _11019_ (.A(_03858_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_03854_),
    .X(_03859_));
 sky130_fd_sc_hd__clkbuf_1 _11021_ (.A(_03859_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_03854_),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_1 _11023_ (.A(_03860_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_03854_),
    .X(_03861_));
 sky130_fd_sc_hd__clkbuf_1 _11025_ (.A(_03861_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_03854_),
    .X(_03862_));
 sky130_fd_sc_hd__clkbuf_1 _11027_ (.A(_03862_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_03854_),
    .X(_03863_));
 sky130_fd_sc_hd__clkbuf_1 _11029_ (.A(_03863_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_03854_),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_1 _11031_ (.A(_03864_),
    .X(_00871_));
 sky130_fd_sc_hd__clkbuf_4 _11032_ (.A(_03717_),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(_03866_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_03865_),
    .X(_03867_));
 sky130_fd_sc_hd__clkbuf_1 _11036_ (.A(_03867_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_03865_),
    .X(_03868_));
 sky130_fd_sc_hd__clkbuf_1 _11038_ (.A(_03868_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_03865_),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_1 _11040_ (.A(_03869_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_03865_),
    .X(_03870_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_03870_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_03865_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_03871_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_03865_),
    .X(_03872_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_03872_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_03865_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_03873_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_03865_),
    .X(_03874_));
 sky130_fd_sc_hd__clkbuf_1 _11050_ (.A(_03874_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_03865_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_1 _11052_ (.A(_03875_),
    .X(_00861_));
 sky130_fd_sc_hd__clkbuf_4 _11053_ (.A(_03717_),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(_03877_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_03876_),
    .X(_03878_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(_03878_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_03876_),
    .X(_03879_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(_03879_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_03876_),
    .X(_03880_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_03880_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_03876_),
    .X(_03881_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_03881_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_03876_),
    .X(_03882_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_03882_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_03876_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_03883_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_03876_),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_03884_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_03876_),
    .X(_03885_));
 sky130_fd_sc_hd__clkbuf_1 _11071_ (.A(_03885_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_03876_),
    .X(_03886_));
 sky130_fd_sc_hd__clkbuf_1 _11073_ (.A(_03886_),
    .X(_00851_));
 sky130_fd_sc_hd__clkbuf_4 _11074_ (.A(_03717_),
    .X(_03887_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(_03888_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_03887_),
    .X(_03889_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(_03889_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_03887_),
    .X(_03890_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(_03890_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_03887_),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_1 _11082_ (.A(_03891_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_03887_),
    .X(_03892_));
 sky130_fd_sc_hd__clkbuf_1 _11084_ (.A(_03892_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_03887_),
    .X(_03893_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(_03893_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_03887_),
    .X(_03894_));
 sky130_fd_sc_hd__clkbuf_1 _11088_ (.A(_03894_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_03887_),
    .X(_03895_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(_03895_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_03887_),
    .X(_03896_));
 sky130_fd_sc_hd__clkbuf_1 _11092_ (.A(_03896_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_03887_),
    .X(_03897_));
 sky130_fd_sc_hd__clkbuf_1 _11094_ (.A(_03897_),
    .X(_00841_));
 sky130_fd_sc_hd__clkbuf_4 _11095_ (.A(_03556_),
    .X(_03898_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_03899_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_03898_),
    .X(_03900_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_03900_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_03898_),
    .X(_03901_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_03901_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_03898_),
    .X(_03902_));
 sky130_fd_sc_hd__clkbuf_1 _11103_ (.A(_03902_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_03898_),
    .X(_03903_));
 sky130_fd_sc_hd__clkbuf_1 _11105_ (.A(_03903_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_03898_),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_1 _11107_ (.A(_03904_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_03898_),
    .X(_03905_));
 sky130_fd_sc_hd__clkbuf_1 _11109_ (.A(_03905_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_03898_),
    .X(_03906_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(_03906_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_03898_),
    .X(_03907_));
 sky130_fd_sc_hd__clkbuf_1 _11113_ (.A(_03907_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _11114_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_03898_),
    .X(_03908_));
 sky130_fd_sc_hd__clkbuf_1 _11115_ (.A(_03908_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_03557_),
    .X(_03909_));
 sky130_fd_sc_hd__clkbuf_1 _11117_ (.A(_03909_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _11118_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_03557_),
    .X(_03910_));
 sky130_fd_sc_hd__clkbuf_1 _11119_ (.A(_03910_),
    .X(_00829_));
 sky130_fd_sc_hd__inv_6 _11120_ (.A(\rbzero.vga_sync.vsync ),
    .Y(net71));
 sky130_fd_sc_hd__buf_6 _11121_ (.A(_03555_),
    .X(_03911_));
 sky130_fd_sc_hd__buf_8 _11122_ (.A(_03911_),
    .X(net60));
 sky130_fd_sc_hd__nand2_4 _11123_ (.A(net71),
    .B(_03480_),
    .Y(_03912_));
 sky130_fd_sc_hd__buf_4 _11124_ (.A(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__buf_4 _11125_ (.A(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__or4_1 _11126_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .B(\rbzero.wall_tracer.visualWallDist[-1] ),
    .C(\rbzero.wall_tracer.visualWallDist[-2] ),
    .D(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_03915_));
 sky130_fd_sc_hd__or4_1 _11127_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(\rbzero.wall_tracer.visualWallDist[7] ),
    .C(\rbzero.wall_tracer.visualWallDist[6] ),
    .D(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_03916_));
 sky130_fd_sc_hd__or4_1 _11128_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(\rbzero.wall_tracer.visualWallDist[3] ),
    .C(\rbzero.wall_tracer.visualWallDist[2] ),
    .D(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_03917_));
 sky130_fd_sc_hd__or4_1 _11129_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(\rbzero.wall_tracer.visualWallDist[9] ),
    .C(_03916_),
    .D(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__clkinv_2 _11130_ (.A(\rbzero.map_rom.f4 ),
    .Y(_03919_));
 sky130_fd_sc_hd__inv_2 _11131_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .Y(_03920_));
 sky130_fd_sc_hd__inv_2 _11132_ (.A(\rbzero.map_rom.a6 ),
    .Y(_03921_));
 sky130_fd_sc_hd__a2bb2o_1 _11133_ (.A1_N(\rbzero.debug_overlay.playerX[0] ),
    .A2_N(_03919_),
    .B1(_03921_),
    .B2(\rbzero.debug_overlay.playerY[3] ),
    .X(_03922_));
 sky130_fd_sc_hd__a221o_1 _11134_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03919_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_03920_),
    .C1(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__clkinv_2 _11135_ (.A(\rbzero.map_rom.f3 ),
    .Y(_03924_));
 sky130_fd_sc_hd__clkinv_2 _11136_ (.A(\rbzero.map_rom.d6 ),
    .Y(_03925_));
 sky130_fd_sc_hd__inv_2 _11137_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .Y(_03926_));
 sky130_fd_sc_hd__a2bb2o_1 _11138_ (.A1_N(\rbzero.debug_overlay.playerY[3] ),
    .A2_N(_03921_),
    .B1(_03926_),
    .B2(\rbzero.map_rom.f3 ),
    .X(_03927_));
 sky130_fd_sc_hd__a221o_1 _11139_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03924_),
    .B1(_03925_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .C1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__clkinv_2 _11140_ (.A(\rbzero.map_rom.f2 ),
    .Y(_03929_));
 sky130_fd_sc_hd__inv_2 _11141_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .Y(_03930_));
 sky130_fd_sc_hd__xor2_1 _11142_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .B(\rbzero.wall_tracer.mapY[5] ),
    .X(_03931_));
 sky130_fd_sc_hd__a221o_1 _11143_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03929_),
    .B1(\rbzero.map_rom.d6 ),
    .B2(_03930_),
    .C1(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__clkbuf_4 _11144_ (.A(\rbzero.map_rom.b6 ),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _11145_ (.A(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__clkinv_2 _11146_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_03935_));
 sky130_fd_sc_hd__clkinv_2 _11147_ (.A(\rbzero.map_rom.f1 ),
    .Y(_03936_));
 sky130_fd_sc_hd__a2bb2o_1 _11148_ (.A1_N(\rbzero.debug_overlay.playerY[2] ),
    .A2_N(_03934_),
    .B1(_03936_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .X(_03937_));
 sky130_fd_sc_hd__a221o_1 _11149_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_03934_),
    .B1(_03935_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .C1(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__or4_2 _11150_ (.A(_03923_),
    .B(_03928_),
    .C(_03932_),
    .D(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__or2_1 _11151_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(\rbzero.wall_tracer.mapX[5] ),
    .X(_03940_));
 sky130_fd_sc_hd__nand2_1 _11152_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(\rbzero.wall_tracer.mapX[5] ),
    .Y(_03941_));
 sky130_fd_sc_hd__buf_2 _11153_ (.A(\rbzero.map_rom.c6 ),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _11154_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__or2_1 _11155_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__xor2_1 _11156_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(\rbzero.map_rom.i_col[4] ),
    .X(_03945_));
 sky130_fd_sc_hd__a221o_1 _11157_ (.A1(_03940_),
    .A2(_03941_),
    .B1(_03943_),
    .B2(_03944_),
    .C1(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__or3_1 _11158_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(\rbzero.wall_tracer.mapX[6] ),
    .C(\rbzero.wall_tracer.mapX[9] ),
    .X(_03947_));
 sky130_fd_sc_hd__o22a_1 _11159_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03929_),
    .B1(_03936_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .X(_03948_));
 sky130_fd_sc_hd__or3b_1 _11160_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_03947_),
    .C_N(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__or4_1 _11161_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(\rbzero.wall_tracer.mapY[8] ),
    .C(\rbzero.wall_tracer.mapY[11] ),
    .D(\rbzero.wall_tracer.mapY[10] ),
    .X(_03950_));
 sky130_fd_sc_hd__or4_1 _11162_ (.A(\rbzero.wall_tracer.mapX[11] ),
    .B(\rbzero.wall_tracer.mapX[10] ),
    .C(\rbzero.wall_tracer.mapY[7] ),
    .D(\rbzero.wall_tracer.mapY[6] ),
    .X(_03951_));
 sky130_fd_sc_hd__or4_1 _11163_ (.A(_03946_),
    .B(_03949_),
    .C(_03950_),
    .D(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__clkinv_4 _11164_ (.A(\rbzero.wall_tracer.visualWallDist[11] ),
    .Y(_03953_));
 sky130_fd_sc_hd__o21a_1 _11165_ (.A1(_03939_),
    .A2(_03952_),
    .B1(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__o21a_1 _11166_ (.A1(_03915_),
    .A2(_03918_),
    .B1(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__xor2_1 _11167_ (.A(\rbzero.otherx[1] ),
    .B(\rbzero.map_rom.f3 ),
    .X(_03956_));
 sky130_fd_sc_hd__a221o_1 _11168_ (.A1(\rbzero.otherx[0] ),
    .A2(_03919_),
    .B1(_03935_),
    .B2(\rbzero.othery[4] ),
    .C1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__inv_2 _11169_ (.A(\rbzero.othery[3] ),
    .Y(_03958_));
 sky130_fd_sc_hd__o2bb2a_1 _11170_ (.A1_N(\rbzero.otherx[2] ),
    .A2_N(_03929_),
    .B1(_03935_),
    .B2(\rbzero.othery[4] ),
    .X(_03959_));
 sky130_fd_sc_hd__o221a_1 _11171_ (.A1(\rbzero.otherx[2] ),
    .A2(_03929_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_03958_),
    .C1(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__xnor2_1 _11172_ (.A(\rbzero.otherx[4] ),
    .B(\rbzero.map_rom.i_col[4] ),
    .Y(_03961_));
 sky130_fd_sc_hd__xnor2_1 _11173_ (.A(\rbzero.othery[2] ),
    .B(_03933_),
    .Y(_03962_));
 sky130_fd_sc_hd__o2bb2a_1 _11174_ (.A1_N(\rbzero.otherx[3] ),
    .A2_N(_03936_),
    .B1(_03919_),
    .B2(\rbzero.otherx[0] ),
    .X(_03963_));
 sky130_fd_sc_hd__o221a_1 _11175_ (.A1(\rbzero.otherx[3] ),
    .A2(_03936_),
    .B1(_03921_),
    .B2(\rbzero.othery[3] ),
    .C1(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__and4_1 _11176_ (.A(_03960_),
    .B(_03961_),
    .C(_03962_),
    .D(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__xnor2_1 _11177_ (.A(\rbzero.othery[0] ),
    .B(\rbzero.map_rom.d6 ),
    .Y(_03966_));
 sky130_fd_sc_hd__xnor2_1 _11178_ (.A(\rbzero.othery[1] ),
    .B(_03942_),
    .Y(_03967_));
 sky130_fd_sc_hd__and4b_2 _11179_ (.A_N(_03957_),
    .B(_03965_),
    .C(_03966_),
    .D(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__and2_1 _11180_ (.A(_03955_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__nand2_1 _11181_ (.A(\rbzero.wall_tracer.state[1] ),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__a22o_1 _11182_ (.A1(\rbzero.map_rom.f3 ),
    .A2(\rbzero.map_rom.f2 ),
    .B1(\rbzero.map_rom.a6 ),
    .B2(\rbzero.map_rom.i_row[4] ),
    .X(_03971_));
 sky130_fd_sc_hd__and4_1 _11183_ (.A(\rbzero.map_rom.d6 ),
    .B(_03942_),
    .C(_03933_),
    .D(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__and3_1 _11184_ (.A(\rbzero.map_rom.f2 ),
    .B(\rbzero.map_rom.f1 ),
    .C(\rbzero.map_rom.i_col[4] ),
    .X(_03973_));
 sky130_fd_sc_hd__nand2_1 _11185_ (.A(\rbzero.map_rom.f2 ),
    .B(_03933_),
    .Y(_03974_));
 sky130_fd_sc_hd__or2_1 _11186_ (.A(\rbzero.map_rom.f2 ),
    .B(_03933_),
    .X(_03975_));
 sky130_fd_sc_hd__nand2_1 _11187_ (.A(_03974_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__or3_1 _11188_ (.A(\rbzero.map_rom.f3 ),
    .B(\rbzero.map_rom.f2 ),
    .C(\rbzero.map_rom.i_col[4] ),
    .X(_03977_));
 sky130_fd_sc_hd__and3b_1 _11189_ (.A_N(_03977_),
    .B(_03936_),
    .C(_03919_),
    .X(_03978_));
 sky130_fd_sc_hd__a31o_1 _11190_ (.A1(_03919_),
    .A2(_03925_),
    .A3(_03976_),
    .B1(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__a31o_1 _11191_ (.A1(\rbzero.map_rom.f4 ),
    .A2(\rbzero.map_rom.f3 ),
    .A3(_03973_),
    .B1(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__o32a_1 _11192_ (.A1(_03933_),
    .A2(\rbzero.map_rom.a6 ),
    .A3(\rbzero.map_rom.i_row[4] ),
    .B1(_03974_),
    .B2(_03924_),
    .X(_03981_));
 sky130_fd_sc_hd__inv_2 _11193_ (.A(_03942_),
    .Y(_03982_));
 sky130_fd_sc_hd__a22o_1 _11194_ (.A1(\rbzero.map_rom.f4 ),
    .A2(\rbzero.map_rom.d6 ),
    .B1(_03982_),
    .B2(_03924_),
    .X(_03983_));
 sky130_fd_sc_hd__a2111o_1 _11195_ (.A1(_03919_),
    .A2(_03925_),
    .B1(\rbzero.map_rom.a6 ),
    .C1(_03983_),
    .D1(\rbzero.map_rom.f1 ),
    .X(_03984_));
 sky130_fd_sc_hd__a211o_1 _11196_ (.A1(\rbzero.map_rom.f3 ),
    .A2(_03942_),
    .B1(_03976_),
    .C1(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__o31a_1 _11197_ (.A1(\rbzero.map_rom.d6 ),
    .A2(_03942_),
    .A3(_03981_),
    .B1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__or3b_4 _11198_ (.A(_03972_),
    .B(_03980_),
    .C_N(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__xnor2_1 _11199_ (.A(\rbzero.map_rom.f4 ),
    .B(_03933_),
    .Y(_03988_));
 sky130_fd_sc_hd__a22o_1 _11200_ (.A1(_03936_),
    .A2(_03982_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(\rbzero.map_rom.f2 ),
    .X(_03989_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(\rbzero.map_rom.f1 ),
    .B(_03942_),
    .Y(_03990_));
 sky130_fd_sc_hd__o22a_1 _11202_ (.A1(_03924_),
    .A2(_03925_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(\rbzero.map_rom.f2 ),
    .X(_03991_));
 sky130_fd_sc_hd__o211a_1 _11203_ (.A1(\rbzero.map_rom.f3 ),
    .A2(\rbzero.map_rom.d6 ),
    .B1(_03990_),
    .C1(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__or3b_1 _11204_ (.A(_03988_),
    .B(_03989_),
    .C_N(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__or4_1 _11205_ (.A(\rbzero.map_rom.f4 ),
    .B(\rbzero.map_rom.d6 ),
    .C(_03921_),
    .D(_03977_),
    .X(_03994_));
 sky130_fd_sc_hd__or4_1 _11206_ (.A(_03933_),
    .B(\rbzero.map_rom.i_row[4] ),
    .C(_03990_),
    .D(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__nand2_2 _11207_ (.A(_03993_),
    .B(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__o21a_1 _11208_ (.A1(_03987_),
    .A2(_03996_),
    .B1(_03955_),
    .X(_03997_));
 sky130_fd_sc_hd__nand2_1 _11209_ (.A(\rbzero.wall_tracer.state[1] ),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__and2_1 _11210_ (.A(_03970_),
    .B(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__nor2_1 _11211_ (.A(_03914_),
    .B(_03999_),
    .Y(_00016_));
 sky130_fd_sc_hd__buf_2 _11212_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_4 _11213_ (.A(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__inv_2 _11214_ (.A(\rbzero.wall_tracer.state[8] ),
    .Y(_04002_));
 sky130_fd_sc_hd__inv_2 _11215_ (.A(\rbzero.wall_tracer.state[11] ),
    .Y(_04003_));
 sky130_fd_sc_hd__a311o_1 _11216_ (.A1(_04001_),
    .A2(_04002_),
    .A3(_04003_),
    .B1(_03914_),
    .C1(\rbzero.wall_tracer.state[0] ),
    .X(_00011_));
 sky130_fd_sc_hd__clkbuf_4 _11217_ (.A(\gpout0.hpos[5] ),
    .X(_04004_));
 sky130_fd_sc_hd__and2_1 _11218_ (.A(\gpout0.hpos[4] ),
    .B(\gpout0.hpos[3] ),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_4 _11219_ (.A(\gpout0.hpos[6] ),
    .X(_04006_));
 sky130_fd_sc_hd__o21ai_1 _11220_ (.A1(_04004_),
    .A2(_04005_),
    .B1(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__and3_1 _11221_ (.A(\gpout0.hpos[5] ),
    .B(\gpout0.hpos[4] ),
    .C(\gpout0.hpos[3] ),
    .X(_04008_));
 sky130_fd_sc_hd__or2_1 _11222_ (.A(\gpout0.hpos[7] ),
    .B(\gpout0.hpos[8] ),
    .X(_04009_));
 sky130_fd_sc_hd__or4b_1 _11223_ (.A(_04007_),
    .B(_04008_),
    .C(_04009_),
    .D_N(_03477_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_4 _11224_ (.A(_04010_),
    .X(net68));
 sky130_fd_sc_hd__inv_2 _11225_ (.A(\gpout0.hpos[7] ),
    .Y(_04011_));
 sky130_fd_sc_hd__a21bo_1 _11226_ (.A1(_04011_),
    .A2(_04007_),
    .B1_N(_03478_),
    .X(net67));
 sky130_fd_sc_hd__inv_2 _11227_ (.A(\rbzero.wall_tracer.state[13] ),
    .Y(_04012_));
 sky130_fd_sc_hd__buf_4 _11228_ (.A(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__buf_4 _11229_ (.A(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__buf_6 _11230_ (.A(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__clkinv_4 _11231_ (.A(\rbzero.wall_tracer.state[1] ),
    .Y(_04016_));
 sky130_fd_sc_hd__or2_2 _11232_ (.A(_04016_),
    .B(_03997_),
    .X(_04017_));
 sky130_fd_sc_hd__or2_1 _11233_ (.A(_03969_),
    .B(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__buf_4 _11234_ (.A(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__a21oi_1 _11235_ (.A1(_04015_),
    .A2(_04019_),
    .B1(_03914_),
    .Y(_00015_));
 sky130_fd_sc_hd__and2_2 _11236_ (.A(\gpout0.hpos[9] ),
    .B(_04009_),
    .X(_04020_));
 sky130_fd_sc_hd__buf_6 _11237_ (.A(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__buf_4 _11238_ (.A(\gpout0.hpos[4] ),
    .X(_04022_));
 sky130_fd_sc_hd__and3_2 _11239_ (.A(\gpout0.hpos[2] ),
    .B(\gpout0.hpos[1] ),
    .C(\gpout0.hpos[0] ),
    .X(_04023_));
 sky130_fd_sc_hd__and2_1 _11240_ (.A(\gpout0.hpos[3] ),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__nor2_1 _11241_ (.A(_03475_),
    .B(_04006_),
    .Y(_04025_));
 sky130_fd_sc_hd__and4b_2 _11242_ (.A_N(_04004_),
    .B(_04022_),
    .C(_04024_),
    .D(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__and3_2 _11243_ (.A(\rbzero.wall_tracer.state[14] ),
    .B(_04021_),
    .C(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_2 _11244_ (.A(_03912_),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__inv_2 _11245_ (.A(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__clkbuf_4 _11246_ (.A(_04029_),
    .X(_00013_));
 sky130_fd_sc_hd__nor2_1 _11247_ (.A(_04003_),
    .B(_03913_),
    .Y(_00000_));
 sky130_fd_sc_hd__buf_2 _11248_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_04030_));
 sky130_fd_sc_hd__buf_2 _11249_ (.A(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__inv_2 _11250_ (.A(\rbzero.wall_tracer.state[0] ),
    .Y(_04032_));
 sky130_fd_sc_hd__nor2_8 _11251_ (.A(\rbzero.vga_sync.vsync ),
    .B(_03555_),
    .Y(_04033_));
 sky130_fd_sc_hd__buf_4 _11252_ (.A(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__buf_4 _11253_ (.A(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__a41o_1 _11254_ (.A1(_04031_),
    .A2(_04032_),
    .A3(_04002_),
    .A4(_04035_),
    .B1(_00000_),
    .X(_00012_));
 sky130_fd_sc_hd__and2_1 _11255_ (.A(_04020_),
    .B(_04026_),
    .X(_04036_));
 sky130_fd_sc_hd__buf_4 _11256_ (.A(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__and2b_1 _11257_ (.A_N(_04037_),
    .B(\rbzero.wall_tracer.state[14] ),
    .X(_04038_));
 sky130_fd_sc_hd__buf_4 _11258_ (.A(_04035_),
    .X(_04039_));
 sky130_fd_sc_hd__o21a_1 _11259_ (.A1(\rbzero.wall_tracer.state[10] ),
    .A2(_04038_),
    .B1(_04039_),
    .X(_00014_));
 sky130_fd_sc_hd__inv_2 _11260_ (.A(\gpout0.vpos[3] ),
    .Y(_04040_));
 sky130_fd_sc_hd__nor2_2 _11261_ (.A(\gpout0.vpos[5] ),
    .B(\gpout0.vpos[4] ),
    .Y(_04041_));
 sky130_fd_sc_hd__nand2_2 _11262_ (.A(_04040_),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__or4_1 _11263_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .D(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__or4b_1 _11264_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(\gpout0.vpos[7] ),
    .D_N(net1),
    .X(_04044_));
 sky130_fd_sc_hd__a21o_1 _11265_ (.A1(_04008_),
    .A2(_04023_),
    .B1(\gpout0.hpos[6] ),
    .X(_04045_));
 sky130_fd_sc_hd__a31oi_4 _11266_ (.A1(\gpout0.hpos[7] ),
    .A2(\gpout0.hpos[8] ),
    .A3(_04045_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04046_));
 sky130_fd_sc_hd__a211o_4 _11267_ (.A1(\gpout0.vpos[6] ),
    .A2(_04043_),
    .B1(_04044_),
    .C1(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__nand2_1 _11268_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_04048_));
 sky130_fd_sc_hd__nand2_1 _11269_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_04049_));
 sky130_fd_sc_hd__or2_1 _11270_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_04050_));
 sky130_fd_sc_hd__nand2_1 _11271_ (.A(_04049_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__or2_1 _11272_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .X(_04052_));
 sky130_fd_sc_hd__nand2_1 _11273_ (.A(_04048_),
    .B(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__or2_1 _11274_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_04054_));
 sky130_fd_sc_hd__nand2_1 _11275_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_04055_));
 sky130_fd_sc_hd__a21boi_1 _11276_ (.A1(\rbzero.texV[8] ),
    .A2(_04054_),
    .B1_N(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__nand2_1 _11277_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_04057_));
 sky130_fd_sc_hd__or2_1 _11278_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_04058_));
 sky130_fd_sc_hd__nand2_1 _11279_ (.A(_04057_),
    .B(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__xor2_1 _11280_ (.A(\rbzero.texV[7] ),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__or2_1 _11281_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_04061_));
 sky130_fd_sc_hd__nand2_1 _11282_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_04062_));
 sky130_fd_sc_hd__a21boi_1 _11283_ (.A1(\rbzero.texV[6] ),
    .A2(_04061_),
    .B1_N(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_1 _11284_ (.A(_04062_),
    .B(_04061_),
    .Y(_04064_));
 sky130_fd_sc_hd__xor2_1 _11285_ (.A(\rbzero.texV[6] ),
    .B(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__or2_1 _11286_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_04066_));
 sky130_fd_sc_hd__nand2_1 _11287_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_04067_));
 sky130_fd_sc_hd__a21boi_1 _11288_ (.A1(\rbzero.texV[5] ),
    .A2(_04066_),
    .B1_N(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2_1 _11289_ (.A(_04065_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand2_1 _11290_ (.A(_04067_),
    .B(_04066_),
    .Y(_04070_));
 sky130_fd_sc_hd__xor2_1 _11291_ (.A(\rbzero.texV[5] ),
    .B(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__or2_1 _11292_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _11293_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_04073_));
 sky130_fd_sc_hd__a21boi_1 _11294_ (.A1(\rbzero.texV[4] ),
    .A2(_04072_),
    .B1_N(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__nor2_1 _11295_ (.A(_04071_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _11296_ (.A(_04073_),
    .B(_04072_),
    .Y(_04076_));
 sky130_fd_sc_hd__xor2_1 _11297_ (.A(\rbzero.texV[4] ),
    .B(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__or2_1 _11298_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_04078_));
 sky130_fd_sc_hd__nand2_1 _11299_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_04079_));
 sky130_fd_sc_hd__a21boi_1 _11300_ (.A1(\rbzero.texV[3] ),
    .A2(_04078_),
    .B1_N(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__nor2_1 _11301_ (.A(_04077_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__xnor2_1 _11302_ (.A(_04077_),
    .B(_04080_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _11303_ (.A(_04079_),
    .B(_04078_),
    .Y(_04083_));
 sky130_fd_sc_hd__xor2_1 _11304_ (.A(\rbzero.texV[3] ),
    .B(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__o211a_1 _11305_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_04085_));
 sky130_fd_sc_hd__a221o_1 _11306_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__o21ai_1 _11307_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__or2_1 _11308_ (.A(_04084_),
    .B(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__nor2_1 _11309_ (.A(_04082_),
    .B(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__and2_1 _11310_ (.A(_04071_),
    .B(_04074_),
    .X(_04090_));
 sky130_fd_sc_hd__or2_1 _11311_ (.A(_04075_),
    .B(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__inv_2 _11312_ (.A(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__o21a_1 _11313_ (.A1(_04081_),
    .A2(_04089_),
    .B1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__and2_1 _11314_ (.A(_04065_),
    .B(_04068_),
    .X(_04094_));
 sky130_fd_sc_hd__or2_1 _11315_ (.A(_04069_),
    .B(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__inv_2 _11316_ (.A(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__o21a_1 _11317_ (.A1(_04075_),
    .A2(_04093_),
    .B1(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__xnor2_1 _11318_ (.A(_04060_),
    .B(_04063_),
    .Y(_04098_));
 sky130_fd_sc_hd__inv_2 _11319_ (.A(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__o21a_1 _11320_ (.A1(_04069_),
    .A2(_04097_),
    .B1(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__o21ba_1 _11321_ (.A1(_04060_),
    .A2(_04063_),
    .B1_N(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__nand2_1 _11322_ (.A(_04055_),
    .B(_04054_),
    .Y(_04102_));
 sky130_fd_sc_hd__xor2_1 _11323_ (.A(\rbzero.texV[8] ),
    .B(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__a21boi_1 _11324_ (.A1(\rbzero.texV[7] ),
    .A2(_04058_),
    .B1_N(_04057_),
    .Y(_04104_));
 sky130_fd_sc_hd__xnor2_1 _11325_ (.A(_04103_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__nor2_1 _11326_ (.A(_04103_),
    .B(_04104_),
    .Y(_04106_));
 sky130_fd_sc_hd__o21ba_1 _11327_ (.A1(_04101_),
    .A2(_04105_),
    .B1_N(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__o21a_1 _11328_ (.A1(_04053_),
    .A2(_04056_),
    .B1(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__a221o_1 _11329_ (.A1(_04048_),
    .A2(_04051_),
    .B1(_04053_),
    .B2(_04056_),
    .C1(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__o21ai_1 _11330_ (.A1(_04048_),
    .A2(_04051_),
    .B1(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__xor2_1 _11331_ (.A(\rbzero.traced_texVinit[11] ),
    .B(\rbzero.texV[11] ),
    .X(_04111_));
 sky130_fd_sc_hd__xnor2_1 _11332_ (.A(_04049_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_2 _11333_ (.A(_04110_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__nor2_8 _11334_ (.A(\rbzero.row_render.vinf ),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__xnor2_1 _11335_ (.A(_04101_),
    .B(_04105_),
    .Y(_04115_));
 sky130_fd_sc_hd__or2_4 _11336_ (.A(_04114_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__nor3_1 _11337_ (.A(_04096_),
    .B(_04075_),
    .C(_04093_),
    .Y(_04117_));
 sky130_fd_sc_hd__or3_1 _11338_ (.A(_04097_),
    .B(_04114_),
    .C(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_4 _11339_ (.A(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__nor3_2 _11340_ (.A(_04099_),
    .B(_04069_),
    .C(_04097_),
    .Y(_04120_));
 sky130_fd_sc_hd__or3_4 _11341_ (.A(_04100_),
    .B(_04114_),
    .C(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__nor3_1 _11342_ (.A(_04092_),
    .B(_04081_),
    .C(_04089_),
    .Y(_04122_));
 sky130_fd_sc_hd__or3_4 _11343_ (.A(_04093_),
    .B(_04114_),
    .C(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__nand2_1 _11344_ (.A(_04082_),
    .B(_04088_),
    .Y(_04124_));
 sky130_fd_sc_hd__or3b_4 _11345_ (.A(_04089_),
    .B(_04114_),
    .C_N(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__buf_4 _11346_ (.A(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__a21oi_1 _11347_ (.A1(_04084_),
    .A2(_04087_),
    .B1(_04114_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _11348_ (.A(_04088_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__buf_4 _11349_ (.A(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__o211a_1 _11350_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04125_),
    .B1(_04129_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_04130_));
 sky130_fd_sc_hd__a221o_1 _11351_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_04123_),
    .B1(_04126_),
    .B2(\rbzero.floor_leak[1] ),
    .C1(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__o221a_1 _11352_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_04123_),
    .B1(_04119_),
    .B2(\rbzero.floor_leak[3] ),
    .C1(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__a221o_1 _11353_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04119_),
    .B1(_04121_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__o22a_1 _11354_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_04121_),
    .B1(_04116_),
    .B2(\rbzero.floor_leak[5] ),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_4 _11355_ (.A(_04088_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_4 _11356_ (.A(_04127_),
    .X(_04136_));
 sky130_fd_sc_hd__and2_1 _11357_ (.A(_04135_),
    .B(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__nor3b_2 _11358_ (.A(_04089_),
    .B(_04114_),
    .C_N(_04124_),
    .Y(_04138_));
 sky130_fd_sc_hd__buf_6 _11359_ (.A(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__clkinv_4 _11360_ (.A(_04116_),
    .Y(_04140_));
 sky130_fd_sc_hd__nor3_2 _11361_ (.A(_04093_),
    .B(_04114_),
    .C(_04122_),
    .Y(_04141_));
 sky130_fd_sc_hd__nor3_4 _11362_ (.A(_04097_),
    .B(_04114_),
    .C(_04117_),
    .Y(_04142_));
 sky130_fd_sc_hd__nor3_4 _11363_ (.A(_04100_),
    .B(_04114_),
    .C(_04120_),
    .Y(_04143_));
 sky130_fd_sc_hd__o21ba_4 _11364_ (.A1(_03476_),
    .A2(_04025_),
    .B1_N(\gpout0.hpos[9] ),
    .X(_04144_));
 sky130_fd_sc_hd__or4_1 _11365_ (.A(_04141_),
    .B(_04142_),
    .C(_04143_),
    .D(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__or4_1 _11366_ (.A(_04137_),
    .B(_04139_),
    .C(_04140_),
    .D(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__inv_2 _11367_ (.A(\rbzero.row_render.size[2] ),
    .Y(_04147_));
 sky130_fd_sc_hd__nor2_1 _11368_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _11369_ (.A(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__or2_1 _11370_ (.A(\rbzero.row_render.size[3] ),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__or3_1 _11371_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__and2_1 _11372_ (.A(\rbzero.row_render.size[6] ),
    .B(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__o21a_1 _11373_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_04152_),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_4 _11374_ (.A(\gpout0.hpos[8] ),
    .X(_04154_));
 sky130_fd_sc_hd__a21o_1 _11375_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04155_));
 sky130_fd_sc_hd__nand3_1 _11376_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .Y(_04156_));
 sky130_fd_sc_hd__and2_1 _11377_ (.A(_04155_),
    .B(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__nor2_1 _11378_ (.A(\rbzero.row_render.size[9] ),
    .B(_04155_),
    .Y(_04158_));
 sky130_fd_sc_hd__xnor2_1 _11379_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_04159_));
 sky130_fd_sc_hd__inv_2 _11380_ (.A(\rbzero.row_render.size[5] ),
    .Y(_04160_));
 sky130_fd_sc_hd__inv_2 _11381_ (.A(\rbzero.row_render.size[4] ),
    .Y(_04161_));
 sky130_fd_sc_hd__inv_2 _11382_ (.A(\rbzero.row_render.size[3] ),
    .Y(_04162_));
 sky130_fd_sc_hd__clkbuf_4 _11383_ (.A(\gpout0.hpos[1] ),
    .X(_04163_));
 sky130_fd_sc_hd__inv_2 _11384_ (.A(\rbzero.row_render.size[1] ),
    .Y(_04164_));
 sky130_fd_sc_hd__inv_2 _11385_ (.A(\rbzero.row_render.size[0] ),
    .Y(_04165_));
 sky130_fd_sc_hd__o211a_1 _11386_ (.A1(_04164_),
    .A2(\gpout0.hpos[1] ),
    .B1(\gpout0.hpos[0] ),
    .C1(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__a221o_1 _11387_ (.A1(_04147_),
    .A2(\gpout0.hpos[2] ),
    .B1(_04163_),
    .B2(_04164_),
    .C1(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__o221a_1 _11388_ (.A1(_04147_),
    .A2(\gpout0.hpos[2] ),
    .B1(\gpout0.hpos[3] ),
    .B2(_04162_),
    .C1(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__a221o_1 _11389_ (.A1(_04161_),
    .A2(_04022_),
    .B1(\gpout0.hpos[3] ),
    .B2(_04162_),
    .C1(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__o221a_1 _11390_ (.A1(_04160_),
    .A2(\gpout0.hpos[5] ),
    .B1(_04022_),
    .B2(_04161_),
    .C1(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__a221o_1 _11391_ (.A1(\rbzero.row_render.size[6] ),
    .A2(\gpout0.hpos[6] ),
    .B1(_04004_),
    .B2(_04160_),
    .C1(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__or2_1 _11392_ (.A(\rbzero.row_render.size[6] ),
    .B(\gpout0.hpos[6] ),
    .X(_04172_));
 sky130_fd_sc_hd__a22o_1 _11393_ (.A1(\gpout0.hpos[7] ),
    .A2(_04159_),
    .B1(_04171_),
    .B2(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__o221a_1 _11394_ (.A1(\gpout0.hpos[7] ),
    .A2(_04159_),
    .B1(_04157_),
    .B2(\gpout0.hpos[8] ),
    .C1(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__a221o_1 _11395_ (.A1(_04154_),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\gpout0.hpos[9] ),
    .C1(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__a21oi_1 _11396_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_04155_),
    .B1(\rbzero.row_render.size[10] ),
    .Y(_04176_));
 sky130_fd_sc_hd__o21a_1 _11397_ (.A1(\gpout0.hpos[9] ),
    .A2(_04158_),
    .B1(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__nor3_1 _11398_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(_04152_),
    .Y(_04178_));
 sky130_fd_sc_hd__nor2_1 _11399_ (.A(_04153_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__nor2_1 _11400_ (.A(\rbzero.row_render.size[9] ),
    .B(_04153_),
    .Y(_04180_));
 sky130_fd_sc_hd__and2_1 _11401_ (.A(\rbzero.row_render.size[9] ),
    .B(_04153_),
    .X(_04181_));
 sky130_fd_sc_hd__xnor2_1 _11402_ (.A(\rbzero.row_render.size[7] ),
    .B(_04152_),
    .Y(_04182_));
 sky130_fd_sc_hd__nor2_1 _11403_ (.A(\rbzero.row_render.size[6] ),
    .B(_04151_),
    .Y(_04183_));
 sky130_fd_sc_hd__nor2_1 _11404_ (.A(_04152_),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__o21ai_1 _11405_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_04150_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_04185_));
 sky130_fd_sc_hd__nand2_1 _11406_ (.A(_04151_),
    .B(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__xnor2_1 _11407_ (.A(\rbzero.row_render.size[4] ),
    .B(_04150_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2_1 _11408_ (.A(\rbzero.row_render.size[3] ),
    .B(_04149_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(_04150_),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__or2_1 _11410_ (.A(_04147_),
    .B(_04148_),
    .X(_04190_));
 sky130_fd_sc_hd__nand3b_1 _11411_ (.A_N(\gpout0.hpos[2] ),
    .B(_04149_),
    .C(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__a21o_1 _11412_ (.A1(\rbzero.row_render.size[0] ),
    .A2(\gpout0.hpos[0] ),
    .B1(_04163_),
    .X(_04192_));
 sky130_fd_sc_hd__a22o_1 _11413_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(_04163_),
    .B2(\gpout0.hpos[0] ),
    .X(_04193_));
 sky130_fd_sc_hd__a211o_1 _11414_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_04192_),
    .B1(_04193_),
    .C1(_04148_),
    .X(_04194_));
 sky130_fd_sc_hd__o211a_1 _11415_ (.A1(\gpout0.hpos[3] ),
    .A2(_04189_),
    .B1(_04191_),
    .C1(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__a221o_1 _11416_ (.A1(\gpout0.hpos[3] ),
    .A2(_04189_),
    .B1(_04187_),
    .B2(_04022_),
    .C1(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__o221a_1 _11417_ (.A1(_04022_),
    .A2(_04187_),
    .B1(_04186_),
    .B2(\gpout0.hpos[5] ),
    .C1(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__a221o_1 _11418_ (.A1(_04004_),
    .A2(_04186_),
    .B1(_04184_),
    .B2(\gpout0.hpos[6] ),
    .C1(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__o221a_1 _11419_ (.A1(\gpout0.hpos[6] ),
    .A2(_04184_),
    .B1(_04182_),
    .B2(\gpout0.hpos[7] ),
    .C1(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__a221o_1 _11420_ (.A1(_03475_),
    .A2(_04182_),
    .B1(_04179_),
    .B2(_04154_),
    .C1(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__o221a_1 _11421_ (.A1(_04154_),
    .A2(_04179_),
    .B1(_04180_),
    .B2(_04181_),
    .C1(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__o2bb2a_1 _11422_ (.A1_N(_04175_),
    .A2_N(_04177_),
    .B1(_04201_),
    .B2(\gpout0.hpos[9] ),
    .X(_04202_));
 sky130_fd_sc_hd__or4_1 _11423_ (.A(\rbzero.row_render.size[10] ),
    .B(\rbzero.row_render.size[9] ),
    .C(_04153_),
    .D(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__a21oi_1 _11424_ (.A1(_04146_),
    .A2(_04203_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04204_));
 sky130_fd_sc_hd__a221o_1 _11425_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_04116_),
    .B1(_04133_),
    .B2(_04134_),
    .C1(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_4 _11426_ (.A(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__buf_6 _11427_ (.A(_04143_),
    .X(_04207_));
 sky130_fd_sc_hd__buf_6 _11428_ (.A(_04141_),
    .X(_04208_));
 sky130_fd_sc_hd__buf_6 _11429_ (.A(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__buf_4 _11430_ (.A(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__buf_4 _11431_ (.A(_04128_),
    .X(_04211_));
 sky130_fd_sc_hd__buf_4 _11432_ (.A(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__buf_4 _11433_ (.A(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_4 _11434_ (.A(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_1 _11435_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__mux2_1 _11436_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04214_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_6 _11437_ (.A(_04125_),
    .X(_04217_));
 sky130_fd_sc_hd__buf_6 _11438_ (.A(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__buf_4 _11439_ (.A(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__mux2_1 _11440_ (.A0(_04215_),
    .A1(_04216_),
    .S(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_4 _11441_ (.A(_04135_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_4 _11442_ (.A(_04136_),
    .X(_04222_));
 sky130_fd_sc_hd__and3_1 _11443_ (.A(\rbzero.tex_r0[57] ),
    .B(_04221_),
    .C(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__buf_4 _11444_ (.A(_04138_),
    .X(_04224_));
 sky130_fd_sc_hd__buf_4 _11445_ (.A(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_4 _11446_ (.A(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__a21o_1 _11447_ (.A1(\rbzero.tex_r0[56] ),
    .A2(_04214_),
    .B1(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__mux2_1 _11448_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04214_),
    .X(_04228_));
 sky130_fd_sc_hd__buf_4 _11449_ (.A(_04123_),
    .X(_04229_));
 sky130_fd_sc_hd__buf_4 _11450_ (.A(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__o221a_1 _11451_ (.A1(_04223_),
    .A2(_04227_),
    .B1(_04228_),
    .B2(_04219_),
    .C1(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__buf_4 _11452_ (.A(_04119_),
    .X(_04232_));
 sky130_fd_sc_hd__a211o_1 _11453_ (.A1(_04210_),
    .A2(_04220_),
    .B1(_04231_),
    .C1(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__mux2_1 _11454_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04214_),
    .X(_04234_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04214_),
    .X(_04235_));
 sky130_fd_sc_hd__mux2_1 _11456_ (.A0(_04234_),
    .A1(_04235_),
    .S(_04226_),
    .X(_04236_));
 sky130_fd_sc_hd__and2_1 _11457_ (.A(\rbzero.tex_r0[54] ),
    .B(_04214_),
    .X(_04237_));
 sky130_fd_sc_hd__a31o_1 _11458_ (.A1(\rbzero.tex_r0[55] ),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04219_),
    .X(_04238_));
 sky130_fd_sc_hd__mux2_1 _11459_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04214_),
    .X(_04239_));
 sky130_fd_sc_hd__o221a_1 _11460_ (.A1(_04237_),
    .A2(_04238_),
    .B1(_04239_),
    .B2(_04226_),
    .C1(_04210_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_8 _11461_ (.A(_04142_),
    .X(_04241_));
 sky130_fd_sc_hd__buf_4 _11462_ (.A(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__a211o_1 _11463_ (.A1(_04230_),
    .A2(_04236_),
    .B1(_04240_),
    .C1(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__buf_4 _11464_ (.A(_04121_),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _11465_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04213_),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04213_),
    .X(_04246_));
 sky130_fd_sc_hd__buf_4 _11467_ (.A(_04139_),
    .X(_04247_));
 sky130_fd_sc_hd__mux2_1 _11468_ (.A0(_04245_),
    .A1(_04246_),
    .S(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__mux2_1 _11469_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04213_),
    .X(_04249_));
 sky130_fd_sc_hd__buf_4 _11470_ (.A(_04211_),
    .X(_04250_));
 sky130_fd_sc_hd__mux2_1 _11471_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__or2_1 _11472_ (.A(_04225_),
    .B(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_8 _11473_ (.A(_04123_),
    .X(_04253_));
 sky130_fd_sc_hd__buf_4 _11474_ (.A(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__o211a_1 _11475_ (.A1(_04219_),
    .A2(_04249_),
    .B1(_04252_),
    .C1(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__a211o_1 _11476_ (.A1(_04210_),
    .A2(_04248_),
    .B1(_04255_),
    .C1(_04232_),
    .X(_04256_));
 sky130_fd_sc_hd__mux2_1 _11477_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04213_),
    .X(_04257_));
 sky130_fd_sc_hd__or2_1 _11478_ (.A(_04226_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04213_),
    .X(_04259_));
 sky130_fd_sc_hd__o21a_1 _11480_ (.A1(_04219_),
    .A2(_04259_),
    .B1(_04254_),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _11481_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04213_),
    .X(_04261_));
 sky130_fd_sc_hd__buf_6 _11482_ (.A(_04211_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_8 _11483_ (.A(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__mux2_1 _11484_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__buf_6 _11485_ (.A(_04126_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_8 _11486_ (.A(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__mux2_1 _11487_ (.A0(_04261_),
    .A1(_04264_),
    .S(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__a221o_1 _11488_ (.A1(_04258_),
    .A2(_04260_),
    .B1(_04267_),
    .B2(_04210_),
    .C1(_04242_),
    .X(_04268_));
 sky130_fd_sc_hd__a31o_1 _11489_ (.A1(_04244_),
    .A2(_04256_),
    .A3(_04268_),
    .B1(_04116_),
    .X(_04269_));
 sky130_fd_sc_hd__a31o_1 _11490_ (.A1(_04207_),
    .A2(_04233_),
    .A3(_04243_),
    .B1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__buf_6 _11491_ (.A(_04129_),
    .X(_04271_));
 sky130_fd_sc_hd__buf_4 _11492_ (.A(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__buf_4 _11493_ (.A(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_1 _11495_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04273_),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _11496_ (.A0(_04274_),
    .A1(_04275_),
    .S(_04226_),
    .X(_04276_));
 sky130_fd_sc_hd__and2_1 _11497_ (.A(\rbzero.tex_r0[14] ),
    .B(_04214_),
    .X(_04277_));
 sky130_fd_sc_hd__a31o_1 _11498_ (.A1(\rbzero.tex_r0[15] ),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04219_),
    .X(_04278_));
 sky130_fd_sc_hd__mux2_1 _11499_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04273_),
    .X(_04279_));
 sky130_fd_sc_hd__o221a_1 _11500_ (.A1(_04277_),
    .A2(_04278_),
    .B1(_04279_),
    .B2(_04226_),
    .C1(_04210_),
    .X(_04280_));
 sky130_fd_sc_hd__a211o_1 _11501_ (.A1(_04230_),
    .A2(_04276_),
    .B1(_04280_),
    .C1(_04232_),
    .X(_04281_));
 sky130_fd_sc_hd__mux2_1 _11502_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04273_),
    .X(_04282_));
 sky130_fd_sc_hd__mux2_1 _11503_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04273_),
    .X(_04283_));
 sky130_fd_sc_hd__mux2_1 _11504_ (.A0(_04282_),
    .A1(_04283_),
    .S(_04226_),
    .X(_04284_));
 sky130_fd_sc_hd__and3_1 _11505_ (.A(\rbzero.tex_r0[3] ),
    .B(_04221_),
    .C(_04222_),
    .X(_04285_));
 sky130_fd_sc_hd__a21o_1 _11506_ (.A1(\rbzero.tex_r0[2] ),
    .A2(_04214_),
    .B1(_04219_),
    .X(_04286_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04273_),
    .X(_04287_));
 sky130_fd_sc_hd__o221a_1 _11508_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04287_),
    .B2(_04226_),
    .C1(_04230_),
    .X(_04288_));
 sky130_fd_sc_hd__a211o_1 _11509_ (.A1(_04210_),
    .A2(_04284_),
    .B1(_04288_),
    .C1(_04242_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_8 _11510_ (.A(_04129_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_8 _11511_ (.A(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__mux2_1 _11512_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04291_),
    .X(_04293_));
 sky130_fd_sc_hd__mux2_1 _11514_ (.A0(_04292_),
    .A1(_04293_),
    .S(_04266_),
    .X(_04294_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04291_),
    .X(_04295_));
 sky130_fd_sc_hd__mux2_1 _11516_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04291_),
    .X(_04296_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(_04295_),
    .A1(_04296_),
    .S(_04247_),
    .X(_04297_));
 sky130_fd_sc_hd__mux2_1 _11518_ (.A0(_04294_),
    .A1(_04297_),
    .S(_04210_),
    .X(_04298_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04263_),
    .X(_04299_));
 sky130_fd_sc_hd__mux2_1 _11520_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04263_),
    .X(_04300_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(_04299_),
    .A1(_04300_),
    .S(_04266_),
    .X(_04301_));
 sky130_fd_sc_hd__mux2_1 _11522_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04213_),
    .X(_04302_));
 sky130_fd_sc_hd__and3_1 _11523_ (.A(\rbzero.tex_r0[31] ),
    .B(_04221_),
    .C(_04222_),
    .X(_04303_));
 sky130_fd_sc_hd__buf_6 _11524_ (.A(_04217_),
    .X(_04304_));
 sky130_fd_sc_hd__a21o_1 _11525_ (.A1(\rbzero.tex_r0[30] ),
    .A2(_04273_),
    .B1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__buf_4 _11526_ (.A(_04209_),
    .X(_04306_));
 sky130_fd_sc_hd__o221a_1 _11527_ (.A1(_04247_),
    .A2(_04302_),
    .B1(_04303_),
    .B2(_04305_),
    .C1(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__a211o_1 _11528_ (.A1(_04230_),
    .A2(_04301_),
    .B1(_04232_),
    .C1(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__o211a_1 _11529_ (.A1(_04242_),
    .A2(_04298_),
    .B1(_04207_),
    .C1(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__a311o_1 _11530_ (.A1(_04244_),
    .A2(_04281_),
    .A3(_04289_),
    .B1(_04309_),
    .C1(_04140_),
    .X(_04310_));
 sky130_fd_sc_hd__nand3b_1 _11531_ (.A_N(_04206_),
    .B(_04270_),
    .C(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__mux2_2 _11532_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_04144_),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _11533_ (.A(_04206_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__clkinv_2 _11534_ (.A(_04047_),
    .Y(_04314_));
 sky130_fd_sc_hd__or2b_4 _11535_ (.A(\gpout0.vpos[5] ),
    .B_N(\gpout0.vpos[4] ),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _11536_ (.A(\gpout0.vpos[5] ),
    .B(\gpout0.vpos[3] ),
    .Y(_04316_));
 sky130_fd_sc_hd__clkbuf_4 _11537_ (.A(\gpout0.hpos[2] ),
    .X(_04317_));
 sky130_fd_sc_hd__and2_1 _11538_ (.A(_04317_),
    .B(_04163_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _11539_ (.A(\gpout0.hpos[0] ),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__o31a_4 _11540_ (.A1(\gpout0.vpos[2] ),
    .A2(\gpout0.vpos[1] ),
    .A3(\gpout0.vpos[0] ),
    .B1(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__o221ai_4 _11541_ (.A1(\gpout0.vpos[3] ),
    .A2(_04315_),
    .B1(_04316_),
    .B2(\gpout0.vpos[4] ),
    .C1(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__and3_1 _11542_ (.A(\gpout0.vpos[8] ),
    .B(\gpout0.vpos[7] ),
    .C(\gpout0.vpos[6] ),
    .X(_04322_));
 sky130_fd_sc_hd__a21o_4 _11543_ (.A1(\gpout0.vpos[5] ),
    .A2(_04322_),
    .B1(\gpout0.vpos[9] ),
    .X(_04323_));
 sky130_fd_sc_hd__a211o_2 _11544_ (.A1(_04314_),
    .A2(_04321_),
    .B1(_04323_),
    .C1(_04020_),
    .X(_04324_));
 sky130_fd_sc_hd__a31o_4 _11545_ (.A1(_04047_),
    .A2(_04311_),
    .A3(_04313_),
    .B1(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__inv_2 _11546_ (.A(_04325_),
    .Y(net65));
 sky130_fd_sc_hd__and2_1 _11547_ (.A(\rbzero.tex_r1[14] ),
    .B(_04213_),
    .X(_04326_));
 sky130_fd_sc_hd__buf_4 _11548_ (.A(_04135_),
    .X(_04327_));
 sky130_fd_sc_hd__buf_4 _11549_ (.A(_04136_),
    .X(_04328_));
 sky130_fd_sc_hd__buf_4 _11550_ (.A(_04126_),
    .X(_04329_));
 sky130_fd_sc_hd__a31o_1 _11551_ (.A1(\rbzero.tex_r1[15] ),
    .A2(_04327_),
    .A3(_04328_),
    .B1(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _11552_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04291_),
    .X(_04331_));
 sky130_fd_sc_hd__buf_4 _11553_ (.A(_04208_),
    .X(_04332_));
 sky130_fd_sc_hd__o221a_1 _11554_ (.A1(_04326_),
    .A2(_04330_),
    .B1(_04331_),
    .B2(_04247_),
    .C1(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__mux2_1 _11555_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04291_),
    .X(_04334_));
 sky130_fd_sc_hd__and3_1 _11556_ (.A(\rbzero.tex_r1[11] ),
    .B(_04327_),
    .C(_04328_),
    .X(_04335_));
 sky130_fd_sc_hd__buf_4 _11557_ (.A(_04128_),
    .X(_04336_));
 sky130_fd_sc_hd__buf_6 _11558_ (.A(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_4 _11559_ (.A(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__a21o_1 _11560_ (.A1(\rbzero.tex_r1[10] ),
    .A2(_04338_),
    .B1(_04304_),
    .X(_04339_));
 sky130_fd_sc_hd__o221a_1 _11561_ (.A1(_04247_),
    .A2(_04334_),
    .B1(_04335_),
    .B2(_04339_),
    .C1(_04254_),
    .X(_04340_));
 sky130_fd_sc_hd__buf_4 _11562_ (.A(_04128_),
    .X(_04341_));
 sky130_fd_sc_hd__buf_6 _11563_ (.A(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _11564_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__mux2_1 _11565_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04342_),
    .X(_04344_));
 sky130_fd_sc_hd__buf_6 _11566_ (.A(_04224_),
    .X(_04345_));
 sky130_fd_sc_hd__mux2_1 _11567_ (.A0(_04343_),
    .A1(_04344_),
    .S(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__buf_4 _11568_ (.A(_04135_),
    .X(_04347_));
 sky130_fd_sc_hd__buf_4 _11569_ (.A(_04136_),
    .X(_04348_));
 sky130_fd_sc_hd__and3_1 _11570_ (.A(\rbzero.tex_r1[3] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_8 _11571_ (.A(_04336_),
    .X(_04350_));
 sky130_fd_sc_hd__a21o_1 _11572_ (.A1(\rbzero.tex_r1[2] ),
    .A2(_04350_),
    .B1(_04217_),
    .X(_04351_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_04342_),
    .X(_04352_));
 sky130_fd_sc_hd__o221a_1 _11574_ (.A1(_04349_),
    .A2(_04351_),
    .B1(_04352_),
    .B2(_04225_),
    .C1(_04253_),
    .X(_04353_));
 sky130_fd_sc_hd__a211o_1 _11575_ (.A1(_04306_),
    .A2(_04346_),
    .B1(_04353_),
    .C1(_04241_),
    .X(_04354_));
 sky130_fd_sc_hd__o311a_1 _11576_ (.A1(_04232_),
    .A2(_04333_),
    .A3(_04340_),
    .B1(_04354_),
    .C1(_04244_),
    .X(_04355_));
 sky130_fd_sc_hd__buf_6 _11577_ (.A(_04341_),
    .X(_04356_));
 sky130_fd_sc_hd__mux2_1 _11578_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__mux2_1 _11579_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04290_),
    .X(_04358_));
 sky130_fd_sc_hd__mux2_1 _11580_ (.A0(_04357_),
    .A1(_04358_),
    .S(_04329_),
    .X(_04359_));
 sky130_fd_sc_hd__mux2_1 _11581_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04290_),
    .X(_04360_));
 sky130_fd_sc_hd__mux2_1 _11582_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04290_),
    .X(_04361_));
 sky130_fd_sc_hd__mux2_1 _11583_ (.A0(_04360_),
    .A1(_04361_),
    .S(_04345_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _11584_ (.A0(_04359_),
    .A1(_04362_),
    .S(_04332_),
    .X(_04363_));
 sky130_fd_sc_hd__mux2_1 _11585_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_04262_),
    .X(_04364_));
 sky130_fd_sc_hd__mux2_1 _11586_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_04342_),
    .X(_04365_));
 sky130_fd_sc_hd__mux2_1 _11587_ (.A0(_04364_),
    .A1(_04365_),
    .S(_04329_),
    .X(_04366_));
 sky130_fd_sc_hd__mux2_1 _11588_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_04342_),
    .X(_04367_));
 sky130_fd_sc_hd__and3_1 _11589_ (.A(\rbzero.tex_r1[31] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04368_));
 sky130_fd_sc_hd__a21o_1 _11590_ (.A1(\rbzero.tex_r1[30] ),
    .A2(_04350_),
    .B1(_04265_),
    .X(_04369_));
 sky130_fd_sc_hd__o221a_1 _11591_ (.A1(_04225_),
    .A2(_04367_),
    .B1(_04368_),
    .B2(_04369_),
    .C1(_04208_),
    .X(_04370_));
 sky130_fd_sc_hd__buf_4 _11592_ (.A(_04119_),
    .X(_04371_));
 sky130_fd_sc_hd__a211o_1 _11593_ (.A1(_04254_),
    .A2(_04366_),
    .B1(_04370_),
    .C1(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__o211a_1 _11594_ (.A1(_04242_),
    .A2(_04363_),
    .B1(_04372_),
    .C1(_04207_),
    .X(_04373_));
 sky130_fd_sc_hd__or3_1 _11595_ (.A(_04140_),
    .B(_04355_),
    .C(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_1 _11596_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_04338_),
    .X(_04375_));
 sky130_fd_sc_hd__mux2_1 _11597_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_04338_),
    .X(_04376_));
 sky130_fd_sc_hd__mux2_1 _11598_ (.A0(_04375_),
    .A1(_04376_),
    .S(_04219_),
    .X(_04377_));
 sky130_fd_sc_hd__and3_1 _11599_ (.A(\rbzero.tex_r1[57] ),
    .B(_04221_),
    .C(_04222_),
    .X(_04378_));
 sky130_fd_sc_hd__buf_4 _11600_ (.A(_04224_),
    .X(_04379_));
 sky130_fd_sc_hd__a21o_1 _11601_ (.A1(\rbzero.tex_r1[56] ),
    .A2(_04273_),
    .B1(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__mux2_1 _11602_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_04338_),
    .X(_04381_));
 sky130_fd_sc_hd__o221a_1 _11603_ (.A1(_04378_),
    .A2(_04380_),
    .B1(_04381_),
    .B2(_04219_),
    .C1(_04230_),
    .X(_04382_));
 sky130_fd_sc_hd__a211o_1 _11604_ (.A1(_04210_),
    .A2(_04377_),
    .B1(_04382_),
    .C1(_04232_),
    .X(_04383_));
 sky130_fd_sc_hd__mux2_1 _11605_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04338_),
    .X(_04384_));
 sky130_fd_sc_hd__mux2_1 _11606_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_04338_),
    .X(_04385_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(_04384_),
    .A1(_04385_),
    .S(_04226_),
    .X(_04386_));
 sky130_fd_sc_hd__and2_1 _11608_ (.A(\rbzero.tex_r1[54] ),
    .B(_04273_),
    .X(_04387_));
 sky130_fd_sc_hd__a31o_1 _11609_ (.A1(\rbzero.tex_r1[55] ),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04266_),
    .X(_04388_));
 sky130_fd_sc_hd__mux2_1 _11610_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_04338_),
    .X(_04389_));
 sky130_fd_sc_hd__o221a_1 _11611_ (.A1(_04387_),
    .A2(_04388_),
    .B1(_04389_),
    .B2(_04226_),
    .C1(_04306_),
    .X(_04390_));
 sky130_fd_sc_hd__a211o_1 _11612_ (.A1(_04230_),
    .A2(_04386_),
    .B1(_04390_),
    .C1(_04242_),
    .X(_04391_));
 sky130_fd_sc_hd__buf_6 _11613_ (.A(_04211_),
    .X(_04392_));
 sky130_fd_sc_hd__mux2_1 _11614_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(_04392_),
    .X(_04394_));
 sky130_fd_sc_hd__mux2_1 _11616_ (.A0(_04393_),
    .A1(_04394_),
    .S(_04304_),
    .X(_04395_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_04392_),
    .X(_04396_));
 sky130_fd_sc_hd__and2_1 _11618_ (.A(\rbzero.tex_r1[46] ),
    .B(_04272_),
    .X(_04397_));
 sky130_fd_sc_hd__a31o_1 _11619_ (.A1(\rbzero.tex_r1[47] ),
    .A2(_04327_),
    .A3(_04328_),
    .B1(_04265_),
    .X(_04398_));
 sky130_fd_sc_hd__o221a_1 _11620_ (.A1(_04379_),
    .A2(_04396_),
    .B1(_04397_),
    .B2(_04398_),
    .C1(_04209_),
    .X(_04399_));
 sky130_fd_sc_hd__a211o_1 _11621_ (.A1(_04230_),
    .A2(_04395_),
    .B1(_04399_),
    .C1(_04371_),
    .X(_04400_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_04392_),
    .X(_04401_));
 sky130_fd_sc_hd__or2_1 _11623_ (.A(_04379_),
    .B(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_1 _11624_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_04350_),
    .X(_04403_));
 sky130_fd_sc_hd__o21a_1 _11625_ (.A1(_04266_),
    .A2(_04403_),
    .B1(_04229_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_1 _11626_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04250_),
    .X(_04405_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_04250_),
    .X(_04406_));
 sky130_fd_sc_hd__mux2_1 _11628_ (.A0(_04405_),
    .A1(_04406_),
    .S(_04218_),
    .X(_04407_));
 sky130_fd_sc_hd__a221o_1 _11629_ (.A1(_04402_),
    .A2(_04404_),
    .B1(_04407_),
    .B2(_04306_),
    .C1(_04241_),
    .X(_04408_));
 sky130_fd_sc_hd__a31o_1 _11630_ (.A1(_04244_),
    .A2(_04400_),
    .A3(_04408_),
    .B1(_04116_),
    .X(_04409_));
 sky130_fd_sc_hd__a31o_1 _11631_ (.A1(_04207_),
    .A2(_04383_),
    .A3(_04391_),
    .B1(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__and3b_1 _11632_ (.A_N(_04206_),
    .B(_04374_),
    .C(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _11633_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_04144_),
    .X(_04412_));
 sky130_fd_sc_hd__a21o_1 _11634_ (.A1(_04206_),
    .A2(_04412_),
    .B1(_04314_),
    .X(_04413_));
 sky130_fd_sc_hd__and3_1 _11635_ (.A(\gpout0.hpos[6] ),
    .B(_04008_),
    .C(_04023_),
    .X(_04414_));
 sky130_fd_sc_hd__a211o_2 _11636_ (.A1(\gpout0.hpos[9] ),
    .A2(_04414_),
    .B1(_04046_),
    .C1(_04020_),
    .X(_04415_));
 sky130_fd_sc_hd__nor2_1 _11637_ (.A(\gpout0.hpos[3] ),
    .B(_04023_),
    .Y(_04416_));
 sky130_fd_sc_hd__or2_2 _11638_ (.A(_04024_),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_1 _11639_ (.A(_04415_),
    .B(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__and2b_1 _11640_ (.A_N(_04022_),
    .B(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__and3b_1 _11641_ (.A_N(_04004_),
    .B(_04419_),
    .C(\gpout0.hpos[6] ),
    .X(_04420_));
 sky130_fd_sc_hd__inv_2 _11642_ (.A(_04414_),
    .Y(_04421_));
 sky130_fd_sc_hd__nand2_4 _11643_ (.A(_04045_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__and2b_1 _11644_ (.A_N(_04415_),
    .B(_04417_),
    .X(_04423_));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__nor2_1 _11646_ (.A(\gpout0.hpos[4] ),
    .B(_04024_),
    .Y(_04425_));
 sky130_fd_sc_hd__a21o_2 _11647_ (.A1(_04005_),
    .A2(_04023_),
    .B1(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__or3_1 _11648_ (.A(\gpout0.hpos[5] ),
    .B(_04424_),
    .C(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__nor2_1 _11649_ (.A(_04422_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__a21oi_1 _11650_ (.A1(_04005_),
    .A2(_04023_),
    .B1(\gpout0.hpos[5] ),
    .Y(_04429_));
 sky130_fd_sc_hd__a21oi_4 _11651_ (.A1(_04008_),
    .A2(_04023_),
    .B1(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__and2_1 _11652_ (.A(_04423_),
    .B(_04426_),
    .X(_04431_));
 sky130_fd_sc_hd__or2b_1 _11653_ (.A(_04430_),
    .B_N(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__nor2_1 _11654_ (.A(_04422_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__and3_1 _11655_ (.A(\gpout0.hpos[6] ),
    .B(_04430_),
    .C(_04431_),
    .X(_04434_));
 sky130_fd_sc_hd__or4_1 _11656_ (.A(_04420_),
    .B(_04428_),
    .C(_04433_),
    .D(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__or4b_2 _11657_ (.A(_04415_),
    .B(_04430_),
    .C(_04417_),
    .D_N(_04022_),
    .X(_04436_));
 sky130_fd_sc_hd__nor2_1 _11658_ (.A(_04422_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_1 _11659_ (.A(_04424_),
    .B(_04426_),
    .Y(_04438_));
 sky130_fd_sc_hd__and2_1 _11660_ (.A(_04004_),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__and2_1 _11661_ (.A(_04418_),
    .B(_04430_),
    .X(_04440_));
 sky130_fd_sc_hd__nor2_1 _11662_ (.A(\gpout0.hpos[7] ),
    .B(_04414_),
    .Y(_04441_));
 sky130_fd_sc_hd__nor2_1 _11663_ (.A(_04011_),
    .B(_04421_),
    .Y(_04442_));
 sky130_fd_sc_hd__nor2_1 _11664_ (.A(_04441_),
    .B(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__and2_2 _11665_ (.A(\gpout0.hpos[8] ),
    .B(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__o41a_1 _11666_ (.A1(_04435_),
    .A2(_04437_),
    .A3(_04439_),
    .A4(_04440_),
    .B1(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__nand2_1 _11667_ (.A(\gpout0.hpos[8] ),
    .B(_04442_),
    .Y(_04446_));
 sky130_fd_sc_hd__a21bo_4 _11668_ (.A1(_03476_),
    .A2(_04441_),
    .B1_N(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__nand2_2 _11669_ (.A(_04422_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__nor2_1 _11670_ (.A(_04427_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__inv_2 _11671_ (.A(_04448_),
    .Y(_04450_));
 sky130_fd_sc_hd__and3b_1 _11672_ (.A_N(_04004_),
    .B(_04419_),
    .C(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__nor2_1 _11673_ (.A(_04432_),
    .B(_04448_),
    .Y(_04452_));
 sky130_fd_sc_hd__or4_4 _11674_ (.A(_04445_),
    .B(_04449_),
    .C(_04451_),
    .D(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__and2_2 _11675_ (.A(_04433_),
    .B(_04447_),
    .X(_04454_));
 sky130_fd_sc_hd__and2_2 _11676_ (.A(_04428_),
    .B(_04447_),
    .X(_04455_));
 sky130_fd_sc_hd__and3_1 _11677_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_04420_),
    .C(_04447_),
    .X(_04456_));
 sky130_fd_sc_hd__a221o_1 _11678_ (.A1(\rbzero.debug_overlay.vplaneX[-5] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .C1(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__and2_2 _11679_ (.A(_04434_),
    .B(_04447_),
    .X(_04458_));
 sky130_fd_sc_hd__nor2_4 _11680_ (.A(_04436_),
    .B(_04448_),
    .Y(_04459_));
 sky130_fd_sc_hd__and3_2 _11681_ (.A(_04004_),
    .B(_04419_),
    .C(_04450_),
    .X(_04460_));
 sky130_fd_sc_hd__a221o_1 _11682_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_04459_),
    .B1(_04460_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .C1(\gpout0.vpos[3] ),
    .X(_04461_));
 sky130_fd_sc_hd__buf_4 _11683_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_04462_));
 sky130_fd_sc_hd__and3_2 _11684_ (.A(_04004_),
    .B(_04438_),
    .C(_04450_),
    .X(_04463_));
 sky130_fd_sc_hd__and3_2 _11685_ (.A(_04022_),
    .B(_04440_),
    .C(_04450_),
    .X(_04464_));
 sky130_fd_sc_hd__and3_2 _11686_ (.A(_04430_),
    .B(_04431_),
    .C(_04450_),
    .X(_04465_));
 sky130_fd_sc_hd__and2_2 _11687_ (.A(_04437_),
    .B(_04447_),
    .X(_04466_));
 sky130_fd_sc_hd__a22o_1 _11688_ (.A1(\rbzero.debug_overlay.vplaneX[-1] ),
    .A2(_04465_),
    .B1(_04466_),
    .B2(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_04467_));
 sky130_fd_sc_hd__a221o_1 _11689_ (.A1(_04462_),
    .A2(_04463_),
    .B1(_04464_),
    .B2(\rbzero.debug_overlay.vplaneX[-4] ),
    .C1(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__a211o_1 _11690_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_04458_),
    .B1(_04461_),
    .C1(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__a211o_1 _11691_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_04453_),
    .B1(_04457_),
    .C1(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__buf_4 _11692_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_04471_));
 sky130_fd_sc_hd__a22o_1 _11693_ (.A1(\rbzero.debug_overlay.vplaneY[-4] ),
    .A2(_04464_),
    .B1(_04460_),
    .B2(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_04472_));
 sky130_fd_sc_hd__a221o_1 _11694_ (.A1(_04471_),
    .A2(_04463_),
    .B1(_04459_),
    .B2(\rbzero.debug_overlay.vplaneY[0] ),
    .C1(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__a221o_1 _11695_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_04455_),
    .B1(_04465_),
    .B2(\rbzero.debug_overlay.vplaneY[-1] ),
    .C1(_04040_),
    .X(_04474_));
 sky130_fd_sc_hd__and2_2 _11696_ (.A(_04420_),
    .B(_04447_),
    .X(_04475_));
 sky130_fd_sc_hd__a22o_1 _11697_ (.A1(\rbzero.debug_overlay.vplaneY[-8] ),
    .A2(_04466_),
    .B1(_04458_),
    .B2(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_04476_));
 sky130_fd_sc_hd__a221o_1 _11698_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(_04475_),
    .B1(_04454_),
    .B2(\rbzero.debug_overlay.vplaneY[-5] ),
    .C1(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__a211o_1 _11699_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_04453_),
    .B1(_04474_),
    .C1(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__o211a_1 _11700_ (.A1(_04473_),
    .A2(_04478_),
    .B1(\gpout0.vpos[5] ),
    .C1(\gpout0.vpos[4] ),
    .X(_04479_));
 sky130_fd_sc_hd__and2_1 _11701_ (.A(_04470_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__or2_1 _11702_ (.A(_04040_),
    .B(_04315_),
    .X(_04481_));
 sky130_fd_sc_hd__a22o_1 _11703_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_04475_),
    .B1(_04458_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .X(_04482_));
 sky130_fd_sc_hd__a22o_1 _11704_ (.A1(\rbzero.debug_overlay.facingY[-4] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .X(_04483_));
 sky130_fd_sc_hd__a22o_1 _11705_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_04459_),
    .B1(_04460_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .X(_04484_));
 sky130_fd_sc_hd__a221o_1 _11706_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_04454_),
    .B1(_04463_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .C1(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__a211o_1 _11707_ (.A1(\rbzero.debug_overlay.facingY[-8] ),
    .A2(_04466_),
    .B1(_04483_),
    .C1(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__a211o_1 _11708_ (.A1(\rbzero.debug_overlay.facingY[-7] ),
    .A2(_04455_),
    .B1(_04482_),
    .C1(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__a21oi_1 _11709_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_04453_),
    .B1(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__or4b_1 _11710_ (.A(\gpout0.vpos[4] ),
    .B(\gpout0.vpos[3] ),
    .C(_04488_),
    .D_N(\gpout0.vpos[5] ),
    .X(_04489_));
 sky130_fd_sc_hd__nand2_1 _11711_ (.A(_04481_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__a22o_1 _11712_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_04464_),
    .B1(_04465_),
    .B2(\rbzero.debug_overlay.facingX[-1] ),
    .X(_04491_));
 sky130_fd_sc_hd__a221o_1 _11713_ (.A1(\rbzero.debug_overlay.facingX[0] ),
    .A2(_04459_),
    .B1(_04460_),
    .B2(\rbzero.debug_overlay.facingX[-2] ),
    .C1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__a221o_1 _11714_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_04463_),
    .B1(_04466_),
    .B2(\rbzero.debug_overlay.facingX[-8] ),
    .C1(_04481_),
    .X(_04493_));
 sky130_fd_sc_hd__a22o_1 _11715_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_04475_),
    .B1(_04458_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .X(_04494_));
 sky130_fd_sc_hd__a221o_1 _11716_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .C1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__a211o_1 _11717_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_04453_),
    .B1(_04493_),
    .C1(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__o22a_1 _11718_ (.A1(_04480_),
    .A2(_04490_),
    .B1(_04492_),
    .B2(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__a22o_1 _11719_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_04454_),
    .B1(_04458_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .X(_04498_));
 sky130_fd_sc_hd__and3_1 _11720_ (.A(_04022_),
    .B(_04444_),
    .C(_04440_),
    .X(_04499_));
 sky130_fd_sc_hd__a22o_1 _11721_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_04449_),
    .B1(_04499_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .X(_04500_));
 sky130_fd_sc_hd__a221o_1 _11722_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_04451_),
    .B1(_04466_),
    .B2(\rbzero.debug_overlay.playerY[-8] ),
    .C1(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__nand2_1 _11723_ (.A(\gpout0.vpos[3] ),
    .B(_04041_),
    .Y(_04502_));
 sky130_fd_sc_hd__a22o_1 _11724_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_04459_),
    .B1(_04460_),
    .B2(\rbzero.debug_overlay.playerY[-2] ),
    .X(_04503_));
 sky130_fd_sc_hd__a211o_1 _11725_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_04463_),
    .B1(_04502_),
    .C1(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__a32o_1 _11726_ (.A1(\rbzero.debug_overlay.playerY[5] ),
    .A2(_04444_),
    .A3(_04439_),
    .B1(_04465_),
    .B2(\rbzero.debug_overlay.playerY[-1] ),
    .X(_04505_));
 sky130_fd_sc_hd__a221o_1 _11727_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_04452_),
    .B1(_04464_),
    .B2(\rbzero.debug_overlay.playerY[-4] ),
    .C1(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__a2111o_1 _11728_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_04455_),
    .B1(_04501_),
    .C1(_04504_),
    .D1(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__a211o_1 _11729_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_04475_),
    .B1(_04498_),
    .C1(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__a22o_1 _11730_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_04475_),
    .B1(_04454_),
    .B2(\rbzero.debug_overlay.playerX[-5] ),
    .X(_04509_));
 sky130_fd_sc_hd__a221o_1 _11731_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_04455_),
    .B1(_04458_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__a22o_1 _11732_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_04449_),
    .B1(_04464_),
    .B2(\rbzero.debug_overlay.playerX[-4] ),
    .X(_04511_));
 sky130_fd_sc_hd__a32o_1 _11733_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_04444_),
    .A3(_04439_),
    .B1(_04452_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .X(_04512_));
 sky130_fd_sc_hd__a221o_1 _11734_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_04466_),
    .B1(_04499_),
    .B2(\rbzero.debug_overlay.playerX[4] ),
    .C1(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__a221o_1 _11735_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_04459_),
    .B1(_04460_),
    .B2(\rbzero.debug_overlay.playerX[-2] ),
    .C1(_04042_),
    .X(_04514_));
 sky130_fd_sc_hd__a221o_1 _11736_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_04451_),
    .B1(_04465_),
    .B2(\rbzero.debug_overlay.playerX[-1] ),
    .C1(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__a2111o_1 _11737_ (.A1(\rbzero.debug_overlay.playerX[-3] ),
    .A2(_04463_),
    .B1(_04511_),
    .C1(_04513_),
    .D1(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__or2_1 _11738_ (.A(_04510_),
    .B(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__and3_1 _11739_ (.A(_04320_),
    .B(_04508_),
    .C(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__o21ai_4 _11740_ (.A1(_04041_),
    .A2(_04497_),
    .B1(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__a21oi_1 _11741_ (.A1(_03478_),
    .A2(_04026_),
    .B1(_04047_),
    .Y(_04520_));
 sky130_fd_sc_hd__a211oi_4 _11742_ (.A1(_04519_),
    .A2(_04520_),
    .B1(_04021_),
    .C1(_04323_),
    .Y(_04521_));
 sky130_fd_sc_hd__o21a_1 _11743_ (.A1(_04411_),
    .A2(_04413_),
    .B1(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__buf_8 _11744_ (.A(_04522_),
    .X(net66));
 sky130_fd_sc_hd__and2_1 _11745_ (.A(\rbzero.tex_g0[14] ),
    .B(_04356_),
    .X(_04523_));
 sky130_fd_sc_hd__a31o_1 _11746_ (.A1(\rbzero.tex_g0[15] ),
    .A2(_04135_),
    .A3(_04136_),
    .B1(_04126_),
    .X(_04524_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04271_),
    .X(_04525_));
 sky130_fd_sc_hd__o221a_1 _11748_ (.A1(_04523_),
    .A2(_04524_),
    .B1(_04525_),
    .B2(_04139_),
    .C1(_04208_),
    .X(_04526_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04271_),
    .X(_04527_));
 sky130_fd_sc_hd__and3_1 _11750_ (.A(\rbzero.tex_g0[11] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04528_));
 sky130_fd_sc_hd__a21o_1 _11751_ (.A1(\rbzero.tex_g0[10] ),
    .A2(_04212_),
    .B1(_04217_),
    .X(_04529_));
 sky130_fd_sc_hd__o221a_1 _11752_ (.A1(_04345_),
    .A2(_04527_),
    .B1(_04528_),
    .B2(_04529_),
    .C1(_04253_),
    .X(_04530_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04129_),
    .X(_04531_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04129_),
    .X(_04532_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(_04531_),
    .A1(_04532_),
    .S(_04138_),
    .X(_04533_));
 sky130_fd_sc_hd__and3_1 _11756_ (.A(\rbzero.tex_g0[3] ),
    .B(_04088_),
    .C(_04127_),
    .X(_04534_));
 sky130_fd_sc_hd__a21o_1 _11757_ (.A1(\rbzero.tex_g0[2] ),
    .A2(_04211_),
    .B1(_04125_),
    .X(_04535_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04341_),
    .X(_04536_));
 sky130_fd_sc_hd__o221a_1 _11759_ (.A1(_04534_),
    .A2(_04535_),
    .B1(_04536_),
    .B2(_04224_),
    .C1(_04123_),
    .X(_04537_));
 sky130_fd_sc_hd__a211o_1 _11760_ (.A1(_04208_),
    .A2(_04533_),
    .B1(_04537_),
    .C1(_04142_),
    .X(_04538_));
 sky130_fd_sc_hd__o311a_1 _11761_ (.A1(_04119_),
    .A2(_04526_),
    .A3(_04530_),
    .B1(_04538_),
    .C1(_04121_),
    .X(_04539_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04129_),
    .X(_04540_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04129_),
    .X(_04541_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(_04540_),
    .A1(_04541_),
    .S(_04126_),
    .X(_04542_));
 sky130_fd_sc_hd__mux2_1 _11765_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04129_),
    .X(_04543_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04129_),
    .X(_04544_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(_04543_),
    .A1(_04544_),
    .S(_04138_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(_04542_),
    .A1(_04545_),
    .S(_04208_),
    .X(_04546_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04341_),
    .X(_04547_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_04341_),
    .X(_04548_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(_04547_),
    .A1(_04548_),
    .S(_04126_),
    .X(_04549_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04129_),
    .X(_04550_));
 sky130_fd_sc_hd__and3_1 _11773_ (.A(\rbzero.tex_g0[31] ),
    .B(_04135_),
    .C(_04136_),
    .X(_04551_));
 sky130_fd_sc_hd__a21o_1 _11774_ (.A1(\rbzero.tex_g0[30] ),
    .A2(_04211_),
    .B1(_04125_),
    .X(_04552_));
 sky130_fd_sc_hd__o221a_1 _11775_ (.A1(_04224_),
    .A2(_04550_),
    .B1(_04551_),
    .B2(_04552_),
    .C1(_04141_),
    .X(_04553_));
 sky130_fd_sc_hd__a211o_1 _11776_ (.A1(_04253_),
    .A2(_04549_),
    .B1(_04553_),
    .C1(_04119_),
    .X(_04554_));
 sky130_fd_sc_hd__o211a_1 _11777_ (.A1(_04142_),
    .A2(_04546_),
    .B1(_04554_),
    .C1(_04143_),
    .X(_04555_));
 sky130_fd_sc_hd__or3_1 _11778_ (.A(_04140_),
    .B(_04539_),
    .C(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__mux2_1 _11779_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04262_),
    .X(_04557_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04262_),
    .X(_04558_));
 sky130_fd_sc_hd__mux2_1 _11781_ (.A0(_04557_),
    .A1(_04558_),
    .S(_04218_),
    .X(_04559_));
 sky130_fd_sc_hd__and3_1 _11782_ (.A(\rbzero.tex_g0[57] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04560_));
 sky130_fd_sc_hd__a21o_1 _11783_ (.A1(\rbzero.tex_g0[56] ),
    .A2(_04350_),
    .B1(_04224_),
    .X(_04561_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04212_),
    .X(_04562_));
 sky130_fd_sc_hd__o221a_1 _11785_ (.A1(_04560_),
    .A2(_04561_),
    .B1(_04562_),
    .B2(_04304_),
    .C1(_04253_),
    .X(_04563_));
 sky130_fd_sc_hd__a211o_1 _11786_ (.A1(_04306_),
    .A2(_04559_),
    .B1(_04563_),
    .C1(_04371_),
    .X(_04564_));
 sky130_fd_sc_hd__mux2_1 _11787_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04262_),
    .X(_04565_));
 sky130_fd_sc_hd__mux2_1 _11788_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04262_),
    .X(_04566_));
 sky130_fd_sc_hd__mux2_1 _11789_ (.A0(_04565_),
    .A1(_04566_),
    .S(_04345_),
    .X(_04567_));
 sky130_fd_sc_hd__and2_1 _11790_ (.A(\rbzero.tex_g0[54] ),
    .B(_04350_),
    .X(_04568_));
 sky130_fd_sc_hd__a31o_1 _11791_ (.A1(\rbzero.tex_g0[55] ),
    .A2(_04347_),
    .A3(_04348_),
    .B1(_04217_),
    .X(_04569_));
 sky130_fd_sc_hd__mux2_1 _11792_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04262_),
    .X(_04570_));
 sky130_fd_sc_hd__o221a_1 _11793_ (.A1(_04568_),
    .A2(_04569_),
    .B1(_04570_),
    .B2(_04225_),
    .C1(_04209_),
    .X(_04571_));
 sky130_fd_sc_hd__a211o_1 _11794_ (.A1(_04254_),
    .A2(_04567_),
    .B1(_04571_),
    .C1(_04241_),
    .X(_04572_));
 sky130_fd_sc_hd__mux2_1 _11795_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04211_),
    .X(_04573_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04341_),
    .X(_04574_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(_04573_),
    .A1(_04574_),
    .S(_04217_),
    .X(_04575_));
 sky130_fd_sc_hd__mux2_1 _11798_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04341_),
    .X(_04576_));
 sky130_fd_sc_hd__and2_1 _11799_ (.A(\rbzero.tex_g0[46] ),
    .B(_04336_),
    .X(_04577_));
 sky130_fd_sc_hd__a31o_1 _11800_ (.A1(\rbzero.tex_g0[47] ),
    .A2(_04135_),
    .A3(_04136_),
    .B1(_04126_),
    .X(_04578_));
 sky130_fd_sc_hd__o221a_1 _11801_ (.A1(_04224_),
    .A2(_04576_),
    .B1(_04577_),
    .B2(_04578_),
    .C1(_04141_),
    .X(_04579_));
 sky130_fd_sc_hd__a211o_1 _11802_ (.A1(_04253_),
    .A2(_04575_),
    .B1(_04579_),
    .C1(_04119_),
    .X(_04580_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04341_),
    .X(_04581_));
 sky130_fd_sc_hd__or2_1 _11804_ (.A(_04224_),
    .B(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__mux2_1 _11805_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04211_),
    .X(_04583_));
 sky130_fd_sc_hd__o21a_1 _11806_ (.A1(_04217_),
    .A2(_04583_),
    .B1(_04123_),
    .X(_04584_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04341_),
    .X(_04585_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04341_),
    .X(_04586_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(_04585_),
    .A1(_04586_),
    .S(_04217_),
    .X(_04587_));
 sky130_fd_sc_hd__a221o_1 _11810_ (.A1(_04582_),
    .A2(_04584_),
    .B1(_04587_),
    .B2(_04208_),
    .C1(_04142_),
    .X(_04588_));
 sky130_fd_sc_hd__a31o_1 _11811_ (.A1(_04121_),
    .A2(_04580_),
    .A3(_04588_),
    .B1(_04116_),
    .X(_04589_));
 sky130_fd_sc_hd__a31o_1 _11812_ (.A1(_04207_),
    .A2(_04564_),
    .A3(_04572_),
    .B1(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__and3b_1 _11813_ (.A_N(_04205_),
    .B(_04556_),
    .C(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__mux2_2 _11814_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_04144_),
    .X(_04592_));
 sky130_fd_sc_hd__a21o_1 _11815_ (.A1(_04206_),
    .A2(_04592_),
    .B1(_04314_),
    .X(_04593_));
 sky130_fd_sc_hd__o21ba_1 _11816_ (.A1(_04591_),
    .A2(_04593_),
    .B1_N(_04324_),
    .X(_04594_));
 sky130_fd_sc_hd__buf_8 _11817_ (.A(_04594_),
    .X(net61));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04212_),
    .X(_04595_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04212_),
    .X(_04596_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(_04595_),
    .A1(_04596_),
    .S(_04345_),
    .X(_04597_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_04212_),
    .X(_04598_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04212_),
    .X(_04599_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(_04598_),
    .A1(_04599_),
    .S(_04218_),
    .X(_04600_));
 sky130_fd_sc_hd__mux2_1 _11824_ (.A0(_04597_),
    .A1(_04600_),
    .S(_04332_),
    .X(_04601_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(\rbzero.tex_g1[63] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04337_),
    .X(_04602_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04392_),
    .X(_04603_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(_04602_),
    .A1(_04603_),
    .S(_04304_),
    .X(_04604_));
 sky130_fd_sc_hd__and3_1 _11828_ (.A(\rbzero.tex_g1[57] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04605_));
 sky130_fd_sc_hd__a21o_1 _11829_ (.A1(\rbzero.tex_g1[56] ),
    .A2(_04272_),
    .B1(_04139_),
    .X(_04606_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_04337_),
    .X(_04607_));
 sky130_fd_sc_hd__o221a_1 _11831_ (.A1(_04605_),
    .A2(_04606_),
    .B1(_04607_),
    .B2(_04266_),
    .C1(_04229_),
    .X(_04608_));
 sky130_fd_sc_hd__a211o_1 _11832_ (.A1(_04306_),
    .A2(_04604_),
    .B1(_04608_),
    .C1(_04371_),
    .X(_04609_));
 sky130_fd_sc_hd__o211a_1 _11833_ (.A1(_04242_),
    .A2(_04601_),
    .B1(_04609_),
    .C1(_04207_),
    .X(_04610_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_04350_),
    .X(_04611_));
 sky130_fd_sc_hd__mux2_1 _11835_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_04350_),
    .X(_04612_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(_04611_),
    .A1(_04612_),
    .S(_04304_),
    .X(_04613_));
 sky130_fd_sc_hd__mux2_1 _11837_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_04337_),
    .X(_04614_));
 sky130_fd_sc_hd__and2_1 _11838_ (.A(\rbzero.tex_g1[46] ),
    .B(_04272_),
    .X(_04615_));
 sky130_fd_sc_hd__a31o_1 _11839_ (.A1(\rbzero.tex_g1[47] ),
    .A2(_04327_),
    .A3(_04328_),
    .B1(_04265_),
    .X(_04616_));
 sky130_fd_sc_hd__o221a_1 _11840_ (.A1(_04379_),
    .A2(_04614_),
    .B1(_04615_),
    .B2(_04616_),
    .C1(_04209_),
    .X(_04617_));
 sky130_fd_sc_hd__a211o_1 _11841_ (.A1(_04230_),
    .A2(_04613_),
    .B1(_04617_),
    .C1(_04232_),
    .X(_04618_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_04337_),
    .X(_04619_));
 sky130_fd_sc_hd__or2_1 _11843_ (.A(_04379_),
    .B(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_04350_),
    .X(_04621_));
 sky130_fd_sc_hd__o21a_1 _11845_ (.A1(_04266_),
    .A2(_04621_),
    .B1(_04229_),
    .X(_04622_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_04392_),
    .X(_04623_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_04392_),
    .X(_04624_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(_04623_),
    .A1(_04624_),
    .S(_04304_),
    .X(_04625_));
 sky130_fd_sc_hd__a221o_1 _11849_ (.A1(_04620_),
    .A2(_04622_),
    .B1(_04625_),
    .B2(_04306_),
    .C1(_04241_),
    .X(_04626_));
 sky130_fd_sc_hd__a31o_1 _11850_ (.A1(_04244_),
    .A2(_04618_),
    .A3(_04626_),
    .B1(_04116_),
    .X(_04627_));
 sky130_fd_sc_hd__nor2_1 _11851_ (.A(_04610_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__and2_1 _11852_ (.A(\rbzero.tex_g1[14] ),
    .B(_04272_),
    .X(_04629_));
 sky130_fd_sc_hd__a31o_1 _11853_ (.A1(\rbzero.tex_g1[15] ),
    .A2(_04327_),
    .A3(_04328_),
    .B1(_04265_),
    .X(_04630_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_04337_),
    .X(_04631_));
 sky130_fd_sc_hd__o221a_1 _11855_ (.A1(_04629_),
    .A2(_04630_),
    .B1(_04631_),
    .B2(_04379_),
    .C1(_04209_),
    .X(_04632_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_04350_),
    .X(_04633_));
 sky130_fd_sc_hd__and3_1 _11857_ (.A(\rbzero.tex_g1[11] ),
    .B(_04327_),
    .C(_04328_),
    .X(_04634_));
 sky130_fd_sc_hd__a21o_1 _11858_ (.A1(\rbzero.tex_g1[10] ),
    .A2(_04291_),
    .B1(_04329_),
    .X(_04635_));
 sky130_fd_sc_hd__o221a_1 _11859_ (.A1(_04379_),
    .A2(_04633_),
    .B1(_04634_),
    .B2(_04635_),
    .C1(_04229_),
    .X(_04636_));
 sky130_fd_sc_hd__mux2_1 _11860_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04336_),
    .X(_04637_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04336_),
    .X(_04638_));
 sky130_fd_sc_hd__mux2_1 _11862_ (.A0(_04637_),
    .A1(_04638_),
    .S(_04224_),
    .X(_04639_));
 sky130_fd_sc_hd__and3_1 _11863_ (.A(\rbzero.tex_g1[3] ),
    .B(_04135_),
    .C(_04136_),
    .X(_04640_));
 sky130_fd_sc_hd__a21o_1 _11864_ (.A1(\rbzero.tex_g1[2] ),
    .A2(_04356_),
    .B1(_04126_),
    .X(_04641_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(_04336_),
    .X(_04642_));
 sky130_fd_sc_hd__o221a_1 _11866_ (.A1(_04640_),
    .A2(_04641_),
    .B1(_04642_),
    .B2(_04139_),
    .C1(_04253_),
    .X(_04643_));
 sky130_fd_sc_hd__a211o_1 _11867_ (.A1(_04209_),
    .A2(_04639_),
    .B1(_04643_),
    .C1(_04142_),
    .X(_04644_));
 sky130_fd_sc_hd__o311a_1 _11868_ (.A1(_04371_),
    .A2(_04632_),
    .A3(_04636_),
    .B1(_04644_),
    .C1(_04244_),
    .X(_04645_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04336_),
    .X(_04646_));
 sky130_fd_sc_hd__mux2_1 _11870_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04211_),
    .X(_04647_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(_04646_),
    .A1(_04647_),
    .S(_04217_),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_1 _11872_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04336_),
    .X(_04649_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04211_),
    .X(_04650_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(_04649_),
    .A1(_04650_),
    .S(_04224_),
    .X(_04651_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(_04648_),
    .A1(_04651_),
    .S(_04209_),
    .X(_04652_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04271_),
    .X(_04653_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04336_),
    .X(_04654_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(_04653_),
    .A1(_04654_),
    .S(_04265_),
    .X(_04655_));
 sky130_fd_sc_hd__mux2_1 _11879_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04336_),
    .X(_04656_));
 sky130_fd_sc_hd__and3_1 _11880_ (.A(\rbzero.tex_g1[31] ),
    .B(_04135_),
    .C(_04136_),
    .X(_04657_));
 sky130_fd_sc_hd__a21o_1 _11881_ (.A1(\rbzero.tex_g1[30] ),
    .A2(_04342_),
    .B1(_04126_),
    .X(_04658_));
 sky130_fd_sc_hd__o221a_1 _11882_ (.A1(_04139_),
    .A2(_04656_),
    .B1(_04657_),
    .B2(_04658_),
    .C1(_04208_),
    .X(_04659_));
 sky130_fd_sc_hd__a211o_1 _11883_ (.A1(_04229_),
    .A2(_04655_),
    .B1(_04659_),
    .C1(_04119_),
    .X(_04660_));
 sky130_fd_sc_hd__o211a_1 _11884_ (.A1(_04241_),
    .A2(_04652_),
    .B1(_04660_),
    .C1(_04143_),
    .X(_04661_));
 sky130_fd_sc_hd__or3_1 _11885_ (.A(_04140_),
    .B(_04645_),
    .C(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__or3b_1 _11886_ (.A(_04628_),
    .B(_04206_),
    .C_N(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__mux2_1 _11887_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_04144_),
    .X(_04664_));
 sky130_fd_sc_hd__a21oi_1 _11888_ (.A1(_04206_),
    .A2(_04664_),
    .B1(_04314_),
    .Y(_04665_));
 sky130_fd_sc_hd__a21bo_4 _11889_ (.A1(_04663_),
    .A2(_04665_),
    .B1_N(_04521_),
    .X(_04666_));
 sky130_fd_sc_hd__clkinv_4 _11890_ (.A(_04666_),
    .Y(net62));
 sky130_fd_sc_hd__and2_1 _11891_ (.A(\rbzero.tex_b0[14] ),
    .B(_04291_),
    .X(_04667_));
 sky130_fd_sc_hd__a31o_1 _11892_ (.A1(\rbzero.tex_b0[15] ),
    .A2(_04327_),
    .A3(_04328_),
    .B1(_04329_),
    .X(_04668_));
 sky130_fd_sc_hd__mux2_1 _11893_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_04272_),
    .X(_04669_));
 sky130_fd_sc_hd__o221a_1 _11894_ (.A1(_04667_),
    .A2(_04668_),
    .B1(_04669_),
    .B2(_04379_),
    .C1(_04332_),
    .X(_04670_));
 sky130_fd_sc_hd__mux2_1 _11895_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04272_),
    .X(_04671_));
 sky130_fd_sc_hd__and3_1 _11896_ (.A(\rbzero.tex_b0[11] ),
    .B(_04327_),
    .C(_04328_),
    .X(_04672_));
 sky130_fd_sc_hd__a21o_1 _11897_ (.A1(\rbzero.tex_b0[10] ),
    .A2(_04213_),
    .B1(_04329_),
    .X(_04673_));
 sky130_fd_sc_hd__o221a_1 _11898_ (.A1(_04247_),
    .A2(_04671_),
    .B1(_04672_),
    .B2(_04673_),
    .C1(_04229_),
    .X(_04674_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04290_),
    .X(_04675_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04290_),
    .X(_04676_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(_04675_),
    .A1(_04676_),
    .S(_04139_),
    .X(_04677_));
 sky130_fd_sc_hd__and3_1 _11902_ (.A(\rbzero.tex_b0[3] ),
    .B(_04135_),
    .C(_04136_),
    .X(_04678_));
 sky130_fd_sc_hd__a21o_1 _11903_ (.A1(\rbzero.tex_b0[2] ),
    .A2(_04262_),
    .B1(_04126_),
    .X(_04679_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04290_),
    .X(_04680_));
 sky130_fd_sc_hd__o221a_1 _11905_ (.A1(_04678_),
    .A2(_04679_),
    .B1(_04680_),
    .B2(_04345_),
    .C1(_04253_),
    .X(_04681_));
 sky130_fd_sc_hd__a211o_1 _11906_ (.A1(_04332_),
    .A2(_04677_),
    .B1(_04681_),
    .C1(_04142_),
    .X(_04682_));
 sky130_fd_sc_hd__o311a_1 _11907_ (.A1(_04232_),
    .A2(_04670_),
    .A3(_04674_),
    .B1(_04682_),
    .C1(_04244_),
    .X(_04683_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_04271_),
    .X(_04684_));
 sky130_fd_sc_hd__mux2_1 _11909_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04271_),
    .X(_04685_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(_04684_),
    .A1(_04685_),
    .S(_04265_),
    .X(_04686_));
 sky130_fd_sc_hd__mux2_1 _11911_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04271_),
    .X(_04687_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_04271_),
    .X(_04688_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(_04687_),
    .A1(_04688_),
    .S(_04139_),
    .X(_04689_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(_04686_),
    .A1(_04689_),
    .S(_04209_),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04290_),
    .X(_04691_));
 sky130_fd_sc_hd__or2_1 _11916_ (.A(_04329_),
    .B(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04290_),
    .X(_04693_));
 sky130_fd_sc_hd__o21a_1 _11918_ (.A1(_04345_),
    .A2(_04693_),
    .B1(_04253_),
    .X(_04694_));
 sky130_fd_sc_hd__mux2_1 _11919_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04271_),
    .X(_04695_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_04271_),
    .X(_04696_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(_04695_),
    .A1(_04696_),
    .S(_04139_),
    .X(_04697_));
 sky130_fd_sc_hd__a221o_1 _11922_ (.A1(_04692_),
    .A2(_04694_),
    .B1(_04697_),
    .B2(_04332_),
    .C1(_04371_),
    .X(_04698_));
 sky130_fd_sc_hd__o211a_1 _11923_ (.A1(_04241_),
    .A2(_04690_),
    .B1(_04698_),
    .C1(_04207_),
    .X(_04699_));
 sky130_fd_sc_hd__or3_1 _11924_ (.A(_04140_),
    .B(_04683_),
    .C(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__mux2_1 _11925_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_04263_),
    .X(_04701_));
 sky130_fd_sc_hd__mux2_1 _11926_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04263_),
    .X(_04702_));
 sky130_fd_sc_hd__mux2_1 _11927_ (.A0(_04701_),
    .A1(_04702_),
    .S(_04266_),
    .X(_04703_));
 sky130_fd_sc_hd__and3_1 _11928_ (.A(\rbzero.tex_b0[57] ),
    .B(_04327_),
    .C(_04328_),
    .X(_04704_));
 sky130_fd_sc_hd__a21o_1 _11929_ (.A1(\rbzero.tex_b0[56] ),
    .A2(_04338_),
    .B1(_04225_),
    .X(_04705_));
 sky130_fd_sc_hd__mux2_1 _11930_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_04263_),
    .X(_04706_));
 sky130_fd_sc_hd__o221a_1 _11931_ (.A1(_04704_),
    .A2(_04705_),
    .B1(_04706_),
    .B2(_04219_),
    .C1(_04254_),
    .X(_04707_));
 sky130_fd_sc_hd__a211o_1 _11932_ (.A1(_04210_),
    .A2(_04703_),
    .B1(_04707_),
    .C1(_04232_),
    .X(_04708_));
 sky130_fd_sc_hd__mux2_1 _11933_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_04263_),
    .X(_04709_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04263_),
    .X(_04710_));
 sky130_fd_sc_hd__mux2_1 _11935_ (.A0(_04709_),
    .A1(_04710_),
    .S(_04247_),
    .X(_04711_));
 sky130_fd_sc_hd__and2_1 _11936_ (.A(\rbzero.tex_b0[54] ),
    .B(_04338_),
    .X(_04712_));
 sky130_fd_sc_hd__a31o_1 _11937_ (.A1(\rbzero.tex_b0[55] ),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04218_),
    .X(_04713_));
 sky130_fd_sc_hd__mux2_1 _11938_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_04263_),
    .X(_04714_));
 sky130_fd_sc_hd__o221a_1 _11939_ (.A1(_04712_),
    .A2(_04713_),
    .B1(_04714_),
    .B2(_04247_),
    .C1(_04306_),
    .X(_04715_));
 sky130_fd_sc_hd__a211o_1 _11940_ (.A1(_04230_),
    .A2(_04711_),
    .B1(_04715_),
    .C1(_04242_),
    .X(_04716_));
 sky130_fd_sc_hd__mux2_1 _11941_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_04342_),
    .X(_04717_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04342_),
    .X(_04718_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(_04717_),
    .A1(_04718_),
    .S(_04329_),
    .X(_04719_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04356_),
    .X(_04720_));
 sky130_fd_sc_hd__and2_1 _11945_ (.A(\rbzero.tex_b0[46] ),
    .B(_04337_),
    .X(_04721_));
 sky130_fd_sc_hd__a31o_1 _11946_ (.A1(\rbzero.tex_b0[47] ),
    .A2(_04347_),
    .A3(_04348_),
    .B1(_04217_),
    .X(_04722_));
 sky130_fd_sc_hd__o221a_1 _11947_ (.A1(_04225_),
    .A2(_04720_),
    .B1(_04721_),
    .B2(_04722_),
    .C1(_04208_),
    .X(_04723_));
 sky130_fd_sc_hd__a211o_1 _11948_ (.A1(_04254_),
    .A2(_04719_),
    .B1(_04723_),
    .C1(_04371_),
    .X(_04724_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_04356_),
    .X(_04725_));
 sky130_fd_sc_hd__or2_1 _11950_ (.A(_04345_),
    .B(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_04262_),
    .X(_04727_));
 sky130_fd_sc_hd__o21a_1 _11952_ (.A1(_04218_),
    .A2(_04727_),
    .B1(_04253_),
    .X(_04728_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_04356_),
    .X(_04729_));
 sky130_fd_sc_hd__mux2_1 _11954_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04356_),
    .X(_04730_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(_04729_),
    .A1(_04730_),
    .S(_04329_),
    .X(_04731_));
 sky130_fd_sc_hd__a221o_1 _11956_ (.A1(_04726_),
    .A2(_04728_),
    .B1(_04731_),
    .B2(_04332_),
    .C1(_04241_),
    .X(_04732_));
 sky130_fd_sc_hd__a31o_1 _11957_ (.A1(_04244_),
    .A2(_04724_),
    .A3(_04732_),
    .B1(_04116_),
    .X(_04733_));
 sky130_fd_sc_hd__a31o_1 _11958_ (.A1(_04207_),
    .A2(_04708_),
    .A3(_04716_),
    .B1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__and3b_1 _11959_ (.A_N(_04206_),
    .B(_04700_),
    .C(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _11960_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_04144_),
    .X(_04736_));
 sky130_fd_sc_hd__a21o_1 _11961_ (.A1(_04206_),
    .A2(_04736_),
    .B1(_04314_),
    .X(_04737_));
 sky130_fd_sc_hd__o21bai_4 _11962_ (.A1(_04735_),
    .A2(_04737_),
    .B1_N(_04324_),
    .Y(_04738_));
 sky130_fd_sc_hd__inv_2 _11963_ (.A(_04738_),
    .Y(net63));
 sky130_fd_sc_hd__mux2_1 _11964_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04356_),
    .X(_04739_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04356_),
    .X(_04740_));
 sky130_fd_sc_hd__mux2_1 _11966_ (.A0(_04739_),
    .A1(_04740_),
    .S(_04329_),
    .X(_04741_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04356_),
    .X(_04742_));
 sky130_fd_sc_hd__mux2_1 _11968_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04290_),
    .X(_04743_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(_04742_),
    .A1(_04743_),
    .S(_04345_),
    .X(_04744_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(_04741_),
    .A1(_04744_),
    .S(_04332_),
    .X(_04745_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04262_),
    .X(_04746_));
 sky130_fd_sc_hd__mux2_1 _11972_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04342_),
    .X(_04747_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(_04746_),
    .A1(_04747_),
    .S(_04218_),
    .X(_04748_));
 sky130_fd_sc_hd__mux2_1 _11974_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04342_),
    .X(_04749_));
 sky130_fd_sc_hd__and3_1 _11975_ (.A(\rbzero.tex_b1[31] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04750_));
 sky130_fd_sc_hd__a21o_1 _11976_ (.A1(\rbzero.tex_b1[30] ),
    .A2(_04272_),
    .B1(_04265_),
    .X(_04751_));
 sky130_fd_sc_hd__o221a_1 _11977_ (.A1(_04225_),
    .A2(_04749_),
    .B1(_04750_),
    .B2(_04751_),
    .C1(_04208_),
    .X(_04752_));
 sky130_fd_sc_hd__a211o_1 _11978_ (.A1(_04254_),
    .A2(_04748_),
    .B1(_04752_),
    .C1(_04371_),
    .X(_04753_));
 sky130_fd_sc_hd__o211a_1 _11979_ (.A1(_04242_),
    .A2(_04745_),
    .B1(_04753_),
    .C1(_04207_),
    .X(_04754_));
 sky130_fd_sc_hd__and2_1 _11980_ (.A(\rbzero.tex_b1[14] ),
    .B(_04338_),
    .X(_04755_));
 sky130_fd_sc_hd__a31o_1 _11981_ (.A1(\rbzero.tex_b1[15] ),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04218_),
    .X(_04756_));
 sky130_fd_sc_hd__mux2_1 _11982_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04291_),
    .X(_04757_));
 sky130_fd_sc_hd__o221a_1 _11983_ (.A1(_04755_),
    .A2(_04756_),
    .B1(_04757_),
    .B2(_04247_),
    .C1(_04332_),
    .X(_04758_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04263_),
    .X(_04759_));
 sky130_fd_sc_hd__and3_1 _11985_ (.A(\rbzero.tex_b1[11] ),
    .B(_04221_),
    .C(_04222_),
    .X(_04760_));
 sky130_fd_sc_hd__a21o_1 _11986_ (.A1(\rbzero.tex_b1[10] ),
    .A2(_04273_),
    .B1(_04304_),
    .X(_04761_));
 sky130_fd_sc_hd__o221a_1 _11987_ (.A1(_04247_),
    .A2(_04759_),
    .B1(_04760_),
    .B2(_04761_),
    .C1(_04254_),
    .X(_04762_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04212_),
    .X(_04763_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04212_),
    .X(_04764_));
 sky130_fd_sc_hd__mux2_1 _11990_ (.A0(_04763_),
    .A1(_04764_),
    .S(_04345_),
    .X(_04765_));
 sky130_fd_sc_hd__and3_1 _11991_ (.A(\rbzero.tex_b1[3] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04766_));
 sky130_fd_sc_hd__a21o_1 _11992_ (.A1(\rbzero.tex_b1[2] ),
    .A2(_04272_),
    .B1(_04265_),
    .X(_04767_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_04250_),
    .X(_04768_));
 sky130_fd_sc_hd__o221a_1 _11994_ (.A1(_04766_),
    .A2(_04767_),
    .B1(_04768_),
    .B2(_04225_),
    .C1(_04229_),
    .X(_04769_));
 sky130_fd_sc_hd__a211o_1 _11995_ (.A1(_04306_),
    .A2(_04765_),
    .B1(_04769_),
    .C1(_04241_),
    .X(_04770_));
 sky130_fd_sc_hd__o311a_1 _11996_ (.A1(_04232_),
    .A2(_04758_),
    .A3(_04762_),
    .B1(_04770_),
    .C1(_04244_),
    .X(_04771_));
 sky130_fd_sc_hd__mux2_1 _11997_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04250_),
    .X(_04772_));
 sky130_fd_sc_hd__mux2_1 _11998_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04250_),
    .X(_04773_));
 sky130_fd_sc_hd__mux2_1 _11999_ (.A0(_04772_),
    .A1(_04773_),
    .S(_04225_),
    .X(_04774_));
 sky130_fd_sc_hd__mux2_1 _12000_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04250_),
    .X(_04775_));
 sky130_fd_sc_hd__mux2_1 _12001_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04212_),
    .X(_04776_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(_04775_),
    .A1(_04776_),
    .S(_04218_),
    .X(_04777_));
 sky130_fd_sc_hd__mux2_1 _12003_ (.A0(_04774_),
    .A1(_04777_),
    .S(_04332_),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04337_),
    .X(_04779_));
 sky130_fd_sc_hd__mux2_1 _12005_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04337_),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(_04779_),
    .A1(_04780_),
    .S(_04304_),
    .X(_04781_));
 sky130_fd_sc_hd__and3_1 _12007_ (.A(\rbzero.tex_b1[57] ),
    .B(_04347_),
    .C(_04348_),
    .X(_04782_));
 sky130_fd_sc_hd__a21o_1 _12008_ (.A1(\rbzero.tex_b1[56] ),
    .A2(_04291_),
    .B1(_04139_),
    .X(_04783_));
 sky130_fd_sc_hd__mux2_1 _12009_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_04350_),
    .X(_04784_));
 sky130_fd_sc_hd__o221a_1 _12010_ (.A1(_04782_),
    .A2(_04783_),
    .B1(_04784_),
    .B2(_04266_),
    .C1(_04229_),
    .X(_04785_));
 sky130_fd_sc_hd__a211o_1 _12011_ (.A1(_04210_),
    .A2(_04781_),
    .B1(_04785_),
    .C1(_04371_),
    .X(_04786_));
 sky130_fd_sc_hd__o211a_1 _12012_ (.A1(_04242_),
    .A2(_04778_),
    .B1(_04786_),
    .C1(_04207_),
    .X(_04787_));
 sky130_fd_sc_hd__mux2_1 _12013_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04392_),
    .X(_04788_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04392_),
    .X(_04789_));
 sky130_fd_sc_hd__mux2_1 _12015_ (.A0(_04788_),
    .A1(_04789_),
    .S(_04304_),
    .X(_04790_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04392_),
    .X(_04791_));
 sky130_fd_sc_hd__and2_1 _12017_ (.A(\rbzero.tex_b1[46] ),
    .B(_04272_),
    .X(_04792_));
 sky130_fd_sc_hd__a31o_1 _12018_ (.A1(\rbzero.tex_b1[47] ),
    .A2(_04327_),
    .A3(_04328_),
    .B1(_04265_),
    .X(_04793_));
 sky130_fd_sc_hd__o221a_1 _12019_ (.A1(_04379_),
    .A2(_04791_),
    .B1(_04792_),
    .B2(_04793_),
    .C1(_04209_),
    .X(_04794_));
 sky130_fd_sc_hd__a211o_1 _12020_ (.A1(_04254_),
    .A2(_04790_),
    .B1(_04794_),
    .C1(_04371_),
    .X(_04795_));
 sky130_fd_sc_hd__mux2_1 _12021_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04250_),
    .X(_04796_));
 sky130_fd_sc_hd__or2_1 _12022_ (.A(_04379_),
    .B(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_04337_),
    .X(_04798_));
 sky130_fd_sc_hd__o21a_1 _12024_ (.A1(_04266_),
    .A2(_04798_),
    .B1(_04229_),
    .X(_04799_));
 sky130_fd_sc_hd__mux2_1 _12025_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04250_),
    .X(_04800_));
 sky130_fd_sc_hd__mux2_1 _12026_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04250_),
    .X(_04801_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(_04800_),
    .A1(_04801_),
    .S(_04218_),
    .X(_04802_));
 sky130_fd_sc_hd__a221o_1 _12028_ (.A1(_04797_),
    .A2(_04799_),
    .B1(_04802_),
    .B2(_04306_),
    .C1(_04241_),
    .X(_04803_));
 sky130_fd_sc_hd__a31o_1 _12029_ (.A1(_04244_),
    .A2(_04795_),
    .A3(_04803_),
    .B1(_04116_),
    .X(_04804_));
 sky130_fd_sc_hd__o32a_1 _12030_ (.A1(_04140_),
    .A2(_04754_),
    .A3(_04771_),
    .B1(_04787_),
    .B2(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__mux2_2 _12031_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_04144_),
    .X(_04806_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(_04805_),
    .A1(_04806_),
    .S(_04206_),
    .X(_04807_));
 sky130_fd_sc_hd__o21a_1 _12033_ (.A1(_04314_),
    .A2(_04807_),
    .B1(_04521_),
    .X(_04808_));
 sky130_fd_sc_hd__buf_8 _12034_ (.A(_04808_),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 _12035_ (.A(\gpout0.hpos[3] ),
    .X(_04809_));
 sky130_fd_sc_hd__nor2_1 _12036_ (.A(_04317_),
    .B(_04163_),
    .Y(_04810_));
 sky130_fd_sc_hd__buf_2 _12037_ (.A(_04004_),
    .X(_04811_));
 sky130_fd_sc_hd__o21ba_1 _12038_ (.A1(_04809_),
    .A2(_04810_),
    .B1_N(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__buf_2 _12039_ (.A(_04022_),
    .X(_04813_));
 sky130_fd_sc_hd__clkbuf_4 _12040_ (.A(_04163_),
    .X(_04814_));
 sky130_fd_sc_hd__or2_1 _12041_ (.A(_04317_),
    .B(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__nor2_1 _12042_ (.A(_04813_),
    .B(_04809_),
    .Y(_04816_));
 sky130_fd_sc_hd__a311o_1 _12043_ (.A1(_04811_),
    .A2(_04813_),
    .A3(_04815_),
    .B1(_04816_),
    .C1(_04005_),
    .X(_04817_));
 sky130_fd_sc_hd__xnor2_2 _12044_ (.A(\rbzero.row_render.wall[0] ),
    .B(\rbzero.row_render.wall[1] ),
    .Y(_04818_));
 sky130_fd_sc_hd__xnor2_1 _12045_ (.A(_04809_),
    .B(_04810_),
    .Y(_04819_));
 sky130_fd_sc_hd__nor2_1 _12046_ (.A(_04318_),
    .B(_04810_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(_04814_),
    .B(_03473_),
    .Y(_04821_));
 sky130_fd_sc_hd__or3b_1 _12048_ (.A(\rbzero.row_render.texu[3] ),
    .B(_03473_),
    .C_N(_04163_),
    .X(_04822_));
 sky130_fd_sc_hd__o21ai_1 _12049_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_04821_),
    .B1(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(\rbzero.row_render.texu[1] ),
    .A1(\rbzero.row_render.texu[0] ),
    .S(_03473_),
    .X(_04824_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(_04814_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(\rbzero.row_render.texu[5] ),
    .A1(\rbzero.row_render.texu[4] ),
    .S(_03473_),
    .X(_04826_));
 sky130_fd_sc_hd__o221ai_1 _12053_ (.A1(\rbzero.row_render.side ),
    .A2(_04821_),
    .B1(_04826_),
    .B2(_04814_),
    .C1(_04820_),
    .Y(_04827_));
 sky130_fd_sc_hd__and3b_1 _12054_ (.A_N(_03473_),
    .B(\rbzero.row_render.wall[0] ),
    .C(_04814_),
    .X(_04828_));
 sky130_fd_sc_hd__o32a_1 _12055_ (.A1(_04820_),
    .A2(_04823_),
    .A3(_04825_),
    .B1(_04827_),
    .B2(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__nor2_1 _12056_ (.A(_04819_),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__a41o_1 _12057_ (.A1(_03474_),
    .A2(_04809_),
    .A3(_04810_),
    .A4(_04818_),
    .B1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__or3b_1 _12058_ (.A(_04812_),
    .B(_04817_),
    .C_N(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__o21ai_1 _12059_ (.A1(_03474_),
    .A2(_04815_),
    .B1(_04005_),
    .Y(_04833_));
 sky130_fd_sc_hd__a21o_1 _12060_ (.A1(_03474_),
    .A2(_04820_),
    .B1(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__a21oi_2 _12061_ (.A1(_04832_),
    .A2(_04834_),
    .B1(net68),
    .Y(net69));
 sky130_fd_sc_hd__buf_1 _12062_ (.A(clknet_opt_5_0_i_clk),
    .X(_04835_));
 sky130_fd_sc_hd__inv_2 _20404__5 (.A(clknet_1_1__leaf__03037_),
    .Y(net126));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(net5),
    .B(net4),
    .X(_04836_));
 sky130_fd_sc_hd__nor2_2 _12065_ (.A(net7),
    .B(net6),
    .Y(_04837_));
 sky130_fd_sc_hd__nor2_2 _12066_ (.A(net3),
    .B(net2),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_1 _12067_ (.A(_04837_),
    .B(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__clkbuf_4 _12068_ (.A(net2),
    .X(_04840_));
 sky130_fd_sc_hd__or2_1 _12069_ (.A(_04840_),
    .B(net61),
    .X(_04841_));
 sky130_fd_sc_hd__nand2_1 _12070_ (.A(_04840_),
    .B(_04666_),
    .Y(_04842_));
 sky130_fd_sc_hd__a31o_1 _12071_ (.A1(net6),
    .A2(_04841_),
    .A3(_04842_),
    .B1(net5),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_1 _12072_ (.A(_04840_),
    .B(_04325_),
    .Y(_04844_));
 sky130_fd_sc_hd__a211o_1 _12073_ (.A1(_04840_),
    .A2(net66),
    .B1(_04844_),
    .C1(net6),
    .X(_04845_));
 sky130_fd_sc_hd__nand2_1 _12074_ (.A(net5),
    .B(net6),
    .Y(_04846_));
 sky130_fd_sc_hd__nor2_1 _12075_ (.A(_04840_),
    .B(_04738_),
    .Y(_04847_));
 sky130_fd_sc_hd__a211o_1 _12076_ (.A1(_04840_),
    .A2(net64),
    .B1(_04846_),
    .C1(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__and4b_1 _12077_ (.A_N(net7),
    .B(_04848_),
    .C(net3),
    .D(net4),
    .X(_04849_));
 sky130_fd_sc_hd__inv_2 _12078_ (.A(net4),
    .Y(_04850_));
 sky130_fd_sc_hd__nor2_1 _12079_ (.A(net5),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__clkinv_2 _12080_ (.A(net2),
    .Y(_04852_));
 sky130_fd_sc_hd__and2_1 _12081_ (.A(net3),
    .B(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__a21o_1 _12082_ (.A1(net51),
    .A2(_04837_),
    .B1(net47),
    .X(_04854_));
 sky130_fd_sc_hd__and2_2 _12083_ (.A(net3),
    .B(net2),
    .X(_04855_));
 sky130_fd_sc_hd__a22o_1 _12084_ (.A1(net46),
    .A2(_04853_),
    .B1(_04854_),
    .B2(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__nor2_2 _12085_ (.A(net3),
    .B(_04852_),
    .Y(_04857_));
 sky130_fd_sc_hd__a22o_1 _12086_ (.A1(net43),
    .A2(_04857_),
    .B1(_04838_),
    .B2(net41),
    .X(_04858_));
 sky130_fd_sc_hd__a22o_1 _12087_ (.A1(net38),
    .A2(_04857_),
    .B1(_04838_),
    .B2(net48),
    .X(_04859_));
 sky130_fd_sc_hd__a221o_1 _12088_ (.A1(net40),
    .A2(_04855_),
    .B1(_04853_),
    .B2(net39),
    .C1(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(_04858_),
    .A1(_04860_),
    .S(net5),
    .X(_04861_));
 sky130_fd_sc_hd__a22o_1 _12090_ (.A1(_04851_),
    .A2(_04856_),
    .B1(_04861_),
    .B2(_04850_),
    .X(_04862_));
 sky130_fd_sc_hd__a22o_1 _12091_ (.A1(net68),
    .A2(_04857_),
    .B1(_04838_),
    .B2(_04323_),
    .X(_04863_));
 sky130_fd_sc_hd__a22o_1 _12092_ (.A1(_04021_),
    .A2(_04855_),
    .B1(_04853_),
    .B2(net42),
    .X(_04864_));
 sky130_fd_sc_hd__nor2_1 _12093_ (.A(net5),
    .B(net4),
    .Y(_04865_));
 sky130_fd_sc_hd__a22o_1 _12094_ (.A1(_04851_),
    .A2(_04863_),
    .B1(_04864_),
    .B2(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__buf_6 _12095_ (.A(net51),
    .X(_04867_));
 sky130_fd_sc_hd__and2_1 _12096_ (.A(_04867_),
    .B(_04837_),
    .X(_04868_));
 sky130_fd_sc_hd__inv_2 _12097_ (.A(net6),
    .Y(_04869_));
 sky130_fd_sc_hd__a32o_1 _12098_ (.A1(_04868_),
    .A2(_04851_),
    .A3(_04855_),
    .B1(_04869_),
    .B2(net7),
    .X(_04870_));
 sky130_fd_sc_hd__o21a_1 _12099_ (.A1(_04862_),
    .A2(_04866_),
    .B1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__a22o_1 _12100_ (.A1(\gpout0.hpos[3] ),
    .A2(_04855_),
    .B1(_04857_),
    .B2(_04163_),
    .X(_04872_));
 sky130_fd_sc_hd__a221o_1 _12101_ (.A1(_04317_),
    .A2(_04853_),
    .B1(_04838_),
    .B2(_03473_),
    .C1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__a31o_1 _12102_ (.A1(net5),
    .A2(net4),
    .A3(_04873_),
    .B1(net6),
    .X(_04874_));
 sky130_fd_sc_hd__mux4_1 _12103_ (.A0(_04813_),
    .A1(_04811_),
    .A2(_04006_),
    .A3(_03475_),
    .S0(net2),
    .S1(net3),
    .X(_04875_));
 sky130_fd_sc_hd__or2_1 _12104_ (.A(net4),
    .B(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__or2_1 _12105_ (.A(net5),
    .B(_04850_),
    .X(_04877_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(_04154_),
    .A1(_03477_),
    .S(_04840_),
    .X(_04878_));
 sky130_fd_sc_hd__a21oi_1 _12107_ (.A1(net3),
    .A2(net4),
    .B1(net5),
    .Y(_04879_));
 sky130_fd_sc_hd__o221a_1 _12108_ (.A1(_04877_),
    .A2(_04878_),
    .B1(_04879_),
    .B2(_04869_),
    .C1(net7),
    .X(_04880_));
 sky130_fd_sc_hd__and3_1 _12109_ (.A(_04874_),
    .B(_04876_),
    .C(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__nor2_1 _12110_ (.A(_04869_),
    .B(_04879_),
    .Y(_04882_));
 sky130_fd_sc_hd__buf_2 _12111_ (.A(\gpout0.vpos[2] ),
    .X(_04883_));
 sky130_fd_sc_hd__buf_2 _12112_ (.A(\gpout0.vpos[3] ),
    .X(_04884_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(_04883_),
    .A1(_04884_),
    .S(_04840_),
    .X(_04885_));
 sky130_fd_sc_hd__buf_2 _12114_ (.A(\gpout0.vpos[6] ),
    .X(_04886_));
 sky130_fd_sc_hd__buf_2 _12115_ (.A(\gpout0.vpos[7] ),
    .X(_04887_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(_04886_),
    .A1(_04887_),
    .S(_04840_),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(\gpout0.vpos[4] ),
    .A1(\gpout0.vpos[5] ),
    .S(_04840_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_4 _12118_ (.A(\gpout0.vpos[9] ),
    .X(_04890_));
 sky130_fd_sc_hd__buf_2 _12119_ (.A(\gpout0.vpos[8] ),
    .X(_04891_));
 sky130_fd_sc_hd__buf_2 _12120_ (.A(\gpout0.vpos[1] ),
    .X(_04892_));
 sky130_fd_sc_hd__mux4_1 _12121_ (.A0(_04890_),
    .A1(_04891_),
    .A2(_04892_),
    .A3(\gpout0.vpos[0] ),
    .S0(_04852_),
    .S1(_04846_),
    .X(_04893_));
 sky130_fd_sc_hd__mux4_2 _12122_ (.A0(_04885_),
    .A1(_04888_),
    .A2(_04889_),
    .A3(_04893_),
    .S0(net4),
    .S1(net3),
    .X(_04894_));
 sky130_fd_sc_hd__and2_1 _12123_ (.A(net49),
    .B(_04838_),
    .X(_04895_));
 sky130_fd_sc_hd__a221o_1 _12124_ (.A1(net52),
    .A2(_04853_),
    .B1(_04857_),
    .B2(net50),
    .C1(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__a221o_2 _12125_ (.A1(_04852_),
    .A2(clknet_1_1__leaf__04835_),
    .B1(_04855_),
    .B2(\gpout0.clk_div[1] ),
    .C1(_04838_),
    .X(_04897_));
 sky130_fd_sc_hd__a21o_2 _12126_ (.A1(_03555_),
    .A2(_04857_),
    .B1(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__a22o_2 _12127_ (.A1(_04851_),
    .A2(_04896_),
    .B1(_04898_),
    .B2(_04865_),
    .X(_04899_));
 sky130_fd_sc_hd__a32o_2 _12128_ (.A1(net7),
    .A2(_04882_),
    .A3(_04894_),
    .B1(_04899_),
    .B2(_04837_),
    .X(_04900_));
 sky130_fd_sc_hd__or3_2 _12129_ (.A(_04871_),
    .B(_04881_),
    .C(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__a31o_2 _12130_ (.A1(_04843_),
    .A2(_04845_),
    .A3(_04849_),
    .B1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__o31a_2 _12131_ (.A1(net61),
    .A2(_04836_),
    .A3(_04839_),
    .B1(_04902_),
    .X(net53));
 sky130_fd_sc_hd__nor2_2 _12132_ (.A(net9),
    .B(net8),
    .Y(_04903_));
 sky130_fd_sc_hd__nor2_2 _12133_ (.A(net12),
    .B(net13),
    .Y(_04904_));
 sky130_fd_sc_hd__nor2_2 _12134_ (.A(net11),
    .B(net10),
    .Y(_04905_));
 sky130_fd_sc_hd__inv_2 _12135_ (.A(net9),
    .Y(_04906_));
 sky130_fd_sc_hd__buf_4 _12136_ (.A(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__clkinv_2 _12137_ (.A(net10),
    .Y(_04908_));
 sky130_fd_sc_hd__inv_2 _12138_ (.A(net8),
    .Y(_04909_));
 sky130_fd_sc_hd__clkbuf_4 _12139_ (.A(net8),
    .X(_04910_));
 sky130_fd_sc_hd__or2_1 _12140_ (.A(_04910_),
    .B(net61),
    .X(_04911_));
 sky130_fd_sc_hd__o211a_1 _12141_ (.A1(_04909_),
    .A2(net62),
    .B1(_04911_),
    .C1(net12),
    .X(_04912_));
 sky130_fd_sc_hd__o211a_1 _12142_ (.A1(_04910_),
    .A2(_04738_),
    .B1(net12),
    .C1(net11),
    .X(_04913_));
 sky130_fd_sc_hd__a21bo_1 _12143_ (.A1(_04910_),
    .A2(net64),
    .B1_N(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__nor2_1 _12144_ (.A(_04910_),
    .B(_04325_),
    .Y(_04915_));
 sky130_fd_sc_hd__a211o_1 _12145_ (.A1(_04910_),
    .A2(net66),
    .B1(_04915_),
    .C1(net12),
    .X(_04916_));
 sky130_fd_sc_hd__o211ai_2 _12146_ (.A1(net11),
    .A2(_04912_),
    .B1(_04914_),
    .C1(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__nor2_4 _12147_ (.A(_04907_),
    .B(net8),
    .Y(_04918_));
 sky130_fd_sc_hd__a22o_1 _12148_ (.A1(net49),
    .A2(_04903_),
    .B1(_04918_),
    .B2(net52),
    .X(_04919_));
 sky130_fd_sc_hd__a31o_1 _12149_ (.A1(net50),
    .A2(_04907_),
    .A3(_04910_),
    .B1(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__and3b_1 _12150_ (.A_N(net11),
    .B(net10),
    .C(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__nor2_1 _12151_ (.A(_04906_),
    .B(_04909_),
    .Y(_04922_));
 sky130_fd_sc_hd__and3_1 _12152_ (.A(\gpout1.clk_div[1] ),
    .B(_04922_),
    .C(_04905_),
    .X(_04923_));
 sky130_fd_sc_hd__and3_2 _12153_ (.A(clknet_1_1__leaf__04835_),
    .B(_04918_),
    .C(_04905_),
    .X(_04924_));
 sky130_fd_sc_hd__a2111o_2 _12154_ (.A1(_04907_),
    .A2(_04905_),
    .B1(_04921_),
    .C1(_04923_),
    .D1(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__a21o_1 _12155_ (.A1(net51),
    .A2(_04904_),
    .B1(net47),
    .X(_04926_));
 sky130_fd_sc_hd__a22o_1 _12156_ (.A1(net46),
    .A2(_04918_),
    .B1(_04922_),
    .B2(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__a31o_1 _12157_ (.A1(_04907_),
    .A2(_04910_),
    .A3(net68),
    .B1(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__a21o_1 _12158_ (.A1(_04323_),
    .A2(_04903_),
    .B1(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__and3b_1 _12159_ (.A_N(net11),
    .B(net10),
    .C(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__inv_2 _12160_ (.A(_04918_),
    .Y(_04931_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(\gpout0.hpos[0] ),
    .A1(_04163_),
    .S(_04910_),
    .X(_04932_));
 sky130_fd_sc_hd__o221a_1 _12162_ (.A1(_04317_),
    .A2(_04931_),
    .B1(_04932_),
    .B2(net9),
    .C1(net11),
    .X(_04933_));
 sky130_fd_sc_hd__o311a_1 _12163_ (.A1(_04809_),
    .A2(_04907_),
    .A3(_04909_),
    .B1(net10),
    .C1(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__and3_1 _12164_ (.A(net38),
    .B(_04907_),
    .C(net8),
    .X(_04935_));
 sky130_fd_sc_hd__a221o_1 _12165_ (.A1(net48),
    .A2(_04903_),
    .B1(_04922_),
    .B2(net40),
    .C1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__a21o_1 _12166_ (.A1(net39),
    .A2(_04918_),
    .B1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(net41),
    .A1(net43),
    .S(net8),
    .X(_04938_));
 sky130_fd_sc_hd__and3_1 _12168_ (.A(_04021_),
    .B(_04922_),
    .C(_04905_),
    .X(_04939_));
 sky130_fd_sc_hd__a31o_1 _12169_ (.A1(_04907_),
    .A2(_04905_),
    .A3(_04938_),
    .B1(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__a311o_1 _12170_ (.A1(net42),
    .A2(_04918_),
    .A3(_04905_),
    .B1(_04940_),
    .C1(net12),
    .X(_04941_));
 sky130_fd_sc_hd__a31o_1 _12171_ (.A1(net11),
    .A2(_04908_),
    .A3(_04937_),
    .B1(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__mux4_1 _12172_ (.A0(_04813_),
    .A1(_04811_),
    .A2(_04006_),
    .A3(_03475_),
    .S0(_04910_),
    .S1(net9),
    .X(_04943_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(_04154_),
    .A1(_03477_),
    .S(net8),
    .X(_04944_));
 sky130_fd_sc_hd__o211a_1 _12174_ (.A1(\gpout0.vpos[0] ),
    .A2(net8),
    .B1(net10),
    .C1(net9),
    .X(_04945_));
 sky130_fd_sc_hd__o21a_1 _12175_ (.A1(_04892_),
    .A2(_04909_),
    .B1(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__a311o_1 _12176_ (.A1(_04907_),
    .A2(net10),
    .A3(_04944_),
    .B1(_04946_),
    .C1(net11),
    .X(_04947_));
 sky130_fd_sc_hd__a21oi_1 _12177_ (.A1(_04908_),
    .A2(_04943_),
    .B1(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__mux4_1 _12178_ (.A0(_04883_),
    .A1(_04884_),
    .A2(\gpout0.vpos[6] ),
    .A3(_04887_),
    .S0(_04910_),
    .S1(net10),
    .X(_04949_));
 sky130_fd_sc_hd__mux4_1 _12179_ (.A0(\gpout0.vpos[4] ),
    .A1(\gpout0.vpos[5] ),
    .A2(_04891_),
    .A3(\gpout0.vpos[9] ),
    .S0(net8),
    .S1(net10),
    .X(_04950_));
 sky130_fd_sc_hd__a21bo_1 _12180_ (.A1(net9),
    .A2(_04950_),
    .B1_N(net11),
    .X(_04951_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(_04907_),
    .A2(_04949_),
    .B1(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__o21ai_1 _12182_ (.A1(_04948_),
    .A2(_04952_),
    .B1(net12),
    .Y(_04953_));
 sky130_fd_sc_hd__and4b_1 _12183_ (.A_N(net11),
    .B(net10),
    .C(_04904_),
    .D(_04867_),
    .X(_04954_));
 sky130_fd_sc_hd__a22o_1 _12184_ (.A1(net13),
    .A2(_04953_),
    .B1(_04954_),
    .B2(_04922_),
    .X(_04955_));
 sky130_fd_sc_hd__o31a_1 _12185_ (.A1(_04930_),
    .A2(_04934_),
    .A3(_04942_),
    .B1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__a21oi_2 _12186_ (.A1(_04904_),
    .A2(_04925_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__o41a_2 _12187_ (.A1(_04907_),
    .A2(_04908_),
    .A3(net13),
    .A4(_04917_),
    .B1(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__a41o_2 _12188_ (.A1(_04666_),
    .A2(_04903_),
    .A3(_04904_),
    .A4(_04905_),
    .B1(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__buf_2 _12190_ (.A(net15),
    .X(_04960_));
 sky130_fd_sc_hd__clkbuf_4 _12191_ (.A(net14),
    .X(_04961_));
 sky130_fd_sc_hd__nor2_1 _12192_ (.A(_04960_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__nor2_1 _12193_ (.A(net17),
    .B(net16),
    .Y(_04963_));
 sky130_fd_sc_hd__nor2_1 _12194_ (.A(net18),
    .B(net19),
    .Y(_04964_));
 sky130_fd_sc_hd__and3_1 _12195_ (.A(_04962_),
    .B(_04963_),
    .C(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__clkbuf_4 _12196_ (.A(_04961_),
    .X(_04966_));
 sky130_fd_sc_hd__nand2_1 _12197_ (.A(_04966_),
    .B(_04666_),
    .Y(_04967_));
 sky130_fd_sc_hd__o211a_1 _12198_ (.A1(_04966_),
    .A2(net61),
    .B1(_04967_),
    .C1(net18),
    .X(_04968_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(net17),
    .B(net18),
    .Y(_04969_));
 sky130_fd_sc_hd__nor2_1 _12200_ (.A(_04966_),
    .B(_04738_),
    .Y(_04970_));
 sky130_fd_sc_hd__a211o_1 _12201_ (.A1(_04966_),
    .A2(net64),
    .B1(_04969_),
    .C1(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(net19),
    .Y(_04972_));
 sky130_fd_sc_hd__nor2_1 _12203_ (.A(_04966_),
    .B(_04325_),
    .Y(_04973_));
 sky130_fd_sc_hd__a211o_1 _12204_ (.A1(_04966_),
    .A2(net66),
    .B1(_04973_),
    .C1(net18),
    .X(_04974_));
 sky130_fd_sc_hd__and4_1 _12205_ (.A(_04960_),
    .B(net16),
    .C(_04972_),
    .D(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__o211a_1 _12206_ (.A1(net17),
    .A2(_04968_),
    .B1(_04971_),
    .C1(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__inv_2 _12207_ (.A(net17),
    .Y(_04977_));
 sky130_fd_sc_hd__and2b_1 _12208_ (.A_N(net15),
    .B(net14),
    .X(_04978_));
 sky130_fd_sc_hd__a22o_1 _12209_ (.A1(_04323_),
    .A2(_04962_),
    .B1(_04978_),
    .B2(net68),
    .X(_04979_));
 sky130_fd_sc_hd__and2b_1 _12210_ (.A_N(_04961_),
    .B(_04960_),
    .X(_04980_));
 sky130_fd_sc_hd__and3_1 _12211_ (.A(_04960_),
    .B(_04961_),
    .C(_04963_),
    .X(_04981_));
 sky130_fd_sc_hd__a32o_1 _12212_ (.A1(net42),
    .A2(_04963_),
    .A3(_04980_),
    .B1(_04981_),
    .B2(_04021_),
    .X(_04982_));
 sky130_fd_sc_hd__a31o_1 _12213_ (.A1(_04977_),
    .A2(net16),
    .A3(_04979_),
    .B1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__and3b_1 _12214_ (.A_N(net18),
    .B(net19),
    .C(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__a21o_1 _12215_ (.A1(_04960_),
    .A2(net16),
    .B1(net17),
    .X(_04985_));
 sky130_fd_sc_hd__nand2_1 _12216_ (.A(net18),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(_04883_),
    .A1(_04884_),
    .S(_04966_),
    .X(_04987_));
 sky130_fd_sc_hd__mux2_1 _12218_ (.A0(_04886_),
    .A1(_04887_),
    .S(_04961_),
    .X(_04988_));
 sky130_fd_sc_hd__buf_2 _12219_ (.A(\gpout0.vpos[4] ),
    .X(_04989_));
 sky130_fd_sc_hd__buf_2 _12220_ (.A(\gpout0.vpos[5] ),
    .X(_04990_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(_04989_),
    .A1(_04990_),
    .S(_04961_),
    .X(_04991_));
 sky130_fd_sc_hd__buf_2 _12222_ (.A(\gpout0.vpos[0] ),
    .X(_04992_));
 sky130_fd_sc_hd__mux4_1 _12223_ (.A0(_04891_),
    .A1(_04992_),
    .A2(_04890_),
    .A3(_04892_),
    .S0(_04969_),
    .S1(_04966_),
    .X(_04993_));
 sky130_fd_sc_hd__mux4_1 _12224_ (.A0(_04987_),
    .A1(_04988_),
    .A2(_04991_),
    .A3(_04993_),
    .S0(net16),
    .S1(_04960_),
    .X(_04994_));
 sky130_fd_sc_hd__and3b_1 _12225_ (.A_N(_04986_),
    .B(_04994_),
    .C(net19),
    .X(_04995_));
 sky130_fd_sc_hd__nand2_1 _12226_ (.A(_04977_),
    .B(net16),
    .Y(_04996_));
 sky130_fd_sc_hd__a22o_1 _12227_ (.A1(net49),
    .A2(_04962_),
    .B1(_04980_),
    .B2(net52),
    .X(_04997_));
 sky130_fd_sc_hd__a21oi_1 _12228_ (.A1(net50),
    .A2(_04978_),
    .B1(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__and3_1 _12229_ (.A(net44),
    .B(_04963_),
    .C(_04978_),
    .X(_04999_));
 sky130_fd_sc_hd__a21oi_1 _12230_ (.A1(\gpout2.clk_div[1] ),
    .A2(_04981_),
    .B1(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__a2111o_2 _12231_ (.A1(net125),
    .A2(_04960_),
    .B1(_04966_),
    .C1(net17),
    .D1(net16),
    .X(_05001_));
 sky130_fd_sc_hd__o211a_2 _12232_ (.A1(_04996_),
    .A2(_04998_),
    .B1(_05000_),
    .C1(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__mux4_1 _12233_ (.A0(_03473_),
    .A1(_04814_),
    .A2(_04317_),
    .A3(_04809_),
    .S0(_04961_),
    .S1(_04960_),
    .X(_05003_));
 sky130_fd_sc_hd__a31o_1 _12234_ (.A1(net17),
    .A2(net16),
    .A3(_05003_),
    .B1(net18),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _12235_ (.A0(_04154_),
    .A1(_03477_),
    .S(_04966_),
    .X(_05005_));
 sky130_fd_sc_hd__mux4_1 _12236_ (.A0(_04813_),
    .A1(_04811_),
    .A2(_04006_),
    .A3(_03475_),
    .S0(_04961_),
    .S1(_04960_),
    .X(_05006_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(net16),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__o2111a_1 _12238_ (.A1(_04996_),
    .A2(_05005_),
    .B1(_04986_),
    .C1(_05007_),
    .D1(net19),
    .X(_05008_));
 sky130_fd_sc_hd__nand2_1 _12239_ (.A(_05004_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand2_1 _12240_ (.A(_04960_),
    .B(_04961_),
    .Y(_05010_));
 sky130_fd_sc_hd__or4b_1 _12241_ (.A(net19),
    .B(_04996_),
    .C(_05010_),
    .D_N(_04867_),
    .X(_05011_));
 sky130_fd_sc_hd__a21oi_1 _12242_ (.A1(_04867_),
    .A2(_04964_),
    .B1(net47),
    .Y(_05012_));
 sky130_fd_sc_hd__o2bb2a_1 _12243_ (.A1_N(net46),
    .A2_N(_04980_),
    .B1(_05012_),
    .B2(_05010_),
    .X(_05013_));
 sky130_fd_sc_hd__mux4_1 _12244_ (.A0(net48),
    .A1(net39),
    .A2(net38),
    .A3(net40),
    .S0(net15),
    .S1(_04961_),
    .X(_05014_));
 sky130_fd_sc_hd__a221o_1 _12245_ (.A1(net41),
    .A2(_04962_),
    .B1(_04978_),
    .B2(net43),
    .C1(net17),
    .X(_05015_));
 sky130_fd_sc_hd__o21ai_1 _12246_ (.A1(_04977_),
    .A2(_05014_),
    .B1(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__o22a_1 _12247_ (.A1(_04996_),
    .A2(_05013_),
    .B1(_05016_),
    .B2(net16),
    .X(_05017_));
 sky130_fd_sc_hd__a211o_1 _12248_ (.A1(_04972_),
    .A2(_05011_),
    .B1(_05017_),
    .C1(net18),
    .X(_05018_));
 sky130_fd_sc_hd__o311a_2 _12249_ (.A1(net18),
    .A2(net19),
    .A3(_05002_),
    .B1(_05009_),
    .C1(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__or3b_2 _12250_ (.A(_04984_),
    .B(_04995_),
    .C_N(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__o2bb2a_2 _12251_ (.A1_N(_04325_),
    .A2_N(_04965_),
    .B1(_04976_),
    .B2(_05020_),
    .X(net55));
 sky130_fd_sc_hd__buf_2 _12252_ (.A(net20),
    .X(_05021_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(_05021_),
    .B(_04666_),
    .Y(_05022_));
 sky130_fd_sc_hd__o211a_1 _12254_ (.A1(_05021_),
    .A2(net61),
    .B1(_05022_),
    .C1(net24),
    .X(_05023_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(net23),
    .B(net24),
    .Y(_05024_));
 sky130_fd_sc_hd__nor2_1 _12256_ (.A(_05021_),
    .B(_04738_),
    .Y(_05025_));
 sky130_fd_sc_hd__a211o_1 _12257_ (.A1(_05021_),
    .A2(net64),
    .B1(_05024_),
    .C1(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__inv_2 _12258_ (.A(net25),
    .Y(_05027_));
 sky130_fd_sc_hd__nor2_1 _12259_ (.A(_05021_),
    .B(_04325_),
    .Y(_05028_));
 sky130_fd_sc_hd__a211o_1 _12260_ (.A1(_05021_),
    .A2(net66),
    .B1(_05028_),
    .C1(net24),
    .X(_05029_));
 sky130_fd_sc_hd__and4_1 _12261_ (.A(net21),
    .B(net22),
    .C(_05027_),
    .D(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__o211a_1 _12262_ (.A1(net23),
    .A2(_05023_),
    .B1(_05026_),
    .C1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__inv_2 _12263_ (.A(net21),
    .Y(_05032_));
 sky130_fd_sc_hd__inv_2 _12264_ (.A(net22),
    .Y(_05033_));
 sky130_fd_sc_hd__inv_2 _12265_ (.A(net24),
    .Y(_05034_));
 sky130_fd_sc_hd__o31a_1 _12266_ (.A1(_05032_),
    .A2(_05033_),
    .A3(_05034_),
    .B1(_05024_),
    .X(_05035_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(_04883_),
    .A1(_04884_),
    .S(_05021_),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_1 _12268_ (.A0(_04886_),
    .A1(_04887_),
    .S(_05021_),
    .X(_05037_));
 sky130_fd_sc_hd__mux2_1 _12269_ (.A0(_04989_),
    .A1(_04990_),
    .S(_05021_),
    .X(_05038_));
 sky130_fd_sc_hd__mux4_1 _12270_ (.A0(_04891_),
    .A1(_04992_),
    .A2(_04890_),
    .A3(_04892_),
    .S0(_05024_),
    .S1(_05021_),
    .X(_05039_));
 sky130_fd_sc_hd__mux4_1 _12271_ (.A0(_05036_),
    .A1(_05037_),
    .A2(_05038_),
    .A3(_05039_),
    .S0(net22),
    .S1(net21),
    .X(_05040_));
 sky130_fd_sc_hd__and3b_1 _12272_ (.A_N(_05035_),
    .B(_05040_),
    .C(net25),
    .X(_05041_));
 sky130_fd_sc_hd__nor2_1 _12273_ (.A(net23),
    .B(_05033_),
    .Y(_05042_));
 sky130_fd_sc_hd__and2_1 _12274_ (.A(_05032_),
    .B(net20),
    .X(_05043_));
 sky130_fd_sc_hd__nor2_2 _12275_ (.A(net21),
    .B(net20),
    .Y(_05044_));
 sky130_fd_sc_hd__a22o_1 _12276_ (.A1(net68),
    .A2(_05043_),
    .B1(_05044_),
    .B2(_04323_),
    .X(_05045_));
 sky130_fd_sc_hd__nor2_2 _12277_ (.A(_05032_),
    .B(net20),
    .Y(_05046_));
 sky130_fd_sc_hd__nor2_1 _12278_ (.A(net23),
    .B(net22),
    .Y(_05047_));
 sky130_fd_sc_hd__and3_1 _12279_ (.A(net42),
    .B(_05046_),
    .C(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__and2_1 _12280_ (.A(net21),
    .B(net20),
    .X(_05049_));
 sky130_fd_sc_hd__and3_1 _12281_ (.A(_04021_),
    .B(_05047_),
    .C(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__a211o_1 _12282_ (.A1(_05042_),
    .A2(_05045_),
    .B1(_05048_),
    .C1(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__and4_1 _12283_ (.A(_04867_),
    .B(_05027_),
    .C(_05042_),
    .D(_05049_),
    .X(_05052_));
 sky130_fd_sc_hd__a31o_1 _12284_ (.A1(_04867_),
    .A2(_05034_),
    .A3(_05027_),
    .B1(net47),
    .X(_05053_));
 sky130_fd_sc_hd__a22o_1 _12285_ (.A1(net46),
    .A2(_05046_),
    .B1(_05049_),
    .B2(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__inv_2 _12286_ (.A(net23),
    .Y(_05055_));
 sky130_fd_sc_hd__a22o_1 _12287_ (.A1(net38),
    .A2(_05043_),
    .B1(_05044_),
    .B2(net48),
    .X(_05056_));
 sky130_fd_sc_hd__a22o_1 _12288_ (.A1(net39),
    .A2(_05046_),
    .B1(_05049_),
    .B2(net40),
    .X(_05057_));
 sky130_fd_sc_hd__a221o_1 _12289_ (.A1(net43),
    .A2(_05043_),
    .B1(_05044_),
    .B2(net41),
    .C1(net23),
    .X(_05058_));
 sky130_fd_sc_hd__o311a_1 _12290_ (.A1(_05055_),
    .A2(_05056_),
    .A3(_05057_),
    .B1(_05058_),
    .C1(_05033_),
    .X(_05059_));
 sky130_fd_sc_hd__a21o_1 _12291_ (.A1(_05042_),
    .A2(_05054_),
    .B1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__o211a_1 _12292_ (.A1(net25),
    .A2(_05052_),
    .B1(_05060_),
    .C1(_05034_),
    .X(_05061_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_05055_),
    .B(net22),
    .Y(_05062_));
 sky130_fd_sc_hd__a22o_1 _12294_ (.A1(net49),
    .A2(_05044_),
    .B1(_05046_),
    .B2(net52),
    .X(_05063_));
 sky130_fd_sc_hd__a21oi_1 _12295_ (.A1(net50),
    .A2(_05043_),
    .B1(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__a22o_1 _12296_ (.A1(net45),
    .A2(_05043_),
    .B1(_05049_),
    .B2(\gpout3.clk_div[1] ),
    .X(_05065_));
 sky130_fd_sc_hd__a2bb2o_1 _12297_ (.A1_N(_05062_),
    .A2_N(_05064_),
    .B1(_05065_),
    .B2(_05047_),
    .X(_05066_));
 sky130_fd_sc_hd__and3_2 _12298_ (.A(clknet_1_1__leaf__04835_),
    .B(_05046_),
    .C(_05047_),
    .X(_05067_));
 sky130_fd_sc_hd__nand2_1 _12299_ (.A(_05044_),
    .B(_05047_),
    .Y(_05068_));
 sky130_fd_sc_hd__or3b_2 _12300_ (.A(_05066_),
    .B(_05067_),
    .C_N(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__a22o_1 _12301_ (.A1(_04163_),
    .A2(_05043_),
    .B1(_05049_),
    .B2(_04809_),
    .X(_05070_));
 sky130_fd_sc_hd__a221o_1 _12302_ (.A1(_03473_),
    .A2(_05044_),
    .B1(_05046_),
    .B2(_04317_),
    .C1(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__a31o_1 _12303_ (.A1(net23),
    .A2(net22),
    .A3(_05071_),
    .B1(net24),
    .X(_05072_));
 sky130_fd_sc_hd__mux4_1 _12304_ (.A0(_04813_),
    .A1(_04811_),
    .A2(_04006_),
    .A3(_03475_),
    .S0(net20),
    .S1(net21),
    .X(_05073_));
 sky130_fd_sc_hd__or2_1 _12305_ (.A(net22),
    .B(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__mux2_1 _12306_ (.A0(_04154_),
    .A1(_03477_),
    .S(net20),
    .X(_05075_));
 sky130_fd_sc_hd__o211a_1 _12307_ (.A1(_05062_),
    .A2(_05075_),
    .B1(_05035_),
    .C1(net25),
    .X(_05076_));
 sky130_fd_sc_hd__and3_1 _12308_ (.A(_05072_),
    .B(_05074_),
    .C(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__a31o_2 _12309_ (.A1(_05034_),
    .A2(_05027_),
    .A3(_05069_),
    .B1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a311o_2 _12310_ (.A1(_05034_),
    .A2(net25),
    .A3(_05051_),
    .B1(_05061_),
    .C1(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__or4_1 _12311_ (.A(net24),
    .B(net25),
    .C(net66),
    .D(_05068_),
    .X(_05080_));
 sky130_fd_sc_hd__o31a_2 _12312_ (.A1(_05031_),
    .A2(_05041_),
    .A3(_05079_),
    .B1(_05080_),
    .X(net56));
 sky130_fd_sc_hd__nor2_1 _12313_ (.A(net30),
    .B(net31),
    .Y(_05081_));
 sky130_fd_sc_hd__clkbuf_4 _12314_ (.A(net27),
    .X(_05082_));
 sky130_fd_sc_hd__clkbuf_4 _12315_ (.A(net26),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_1 _12316_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__nor2_1 _12317_ (.A(net29),
    .B(net28),
    .Y(_05085_));
 sky130_fd_sc_hd__and3_1 _12318_ (.A(_05081_),
    .B(_05084_),
    .C(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_4 _12319_ (.A(_05083_),
    .X(_05087_));
 sky130_fd_sc_hd__nand2_1 _12320_ (.A(_05087_),
    .B(_04666_),
    .Y(_05088_));
 sky130_fd_sc_hd__o211a_1 _12321_ (.A1(_05087_),
    .A2(net61),
    .B1(_05088_),
    .C1(net30),
    .X(_05089_));
 sky130_fd_sc_hd__inv_2 _12322_ (.A(net31),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2_1 _12323_ (.A(net29),
    .B(net30),
    .Y(_05091_));
 sky130_fd_sc_hd__nor2_1 _12324_ (.A(_05087_),
    .B(_04738_),
    .Y(_05092_));
 sky130_fd_sc_hd__a211o_1 _12325_ (.A1(_05087_),
    .A2(net64),
    .B1(_05091_),
    .C1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__and2_1 _12326_ (.A(_05082_),
    .B(net28),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _12327_ (.A(_05087_),
    .B(_04325_),
    .Y(_05095_));
 sky130_fd_sc_hd__a211o_1 _12328_ (.A1(_05087_),
    .A2(net66),
    .B1(_05095_),
    .C1(net30),
    .X(_05096_));
 sky130_fd_sc_hd__and4_1 _12329_ (.A(_05090_),
    .B(_05093_),
    .C(_05094_),
    .D(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__o21a_1 _12330_ (.A1(net29),
    .A2(_05089_),
    .B1(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__nand2_1 _12331_ (.A(_05082_),
    .B(_05087_),
    .Y(_05099_));
 sky130_fd_sc_hd__inv_2 _12332_ (.A(net29),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _12333_ (.A(_05100_),
    .B(net28),
    .Y(_05101_));
 sky130_fd_sc_hd__or4b_1 _12334_ (.A(net31),
    .B(_05099_),
    .C(_05101_),
    .D_N(_04867_),
    .X(_05102_));
 sky130_fd_sc_hd__and2b_1 _12335_ (.A_N(_05083_),
    .B(_05082_),
    .X(_05103_));
 sky130_fd_sc_hd__a21oi_1 _12336_ (.A1(_04867_),
    .A2(_05081_),
    .B1(net47),
    .Y(_05104_));
 sky130_fd_sc_hd__o2bb2a_1 _12337_ (.A1_N(net46),
    .A2_N(_05103_),
    .B1(_05104_),
    .B2(_05099_),
    .X(_05105_));
 sky130_fd_sc_hd__mux4_1 _12338_ (.A0(net48),
    .A1(net39),
    .A2(net38),
    .A3(net40),
    .S0(_05082_),
    .S1(_05087_),
    .X(_05106_));
 sky130_fd_sc_hd__and2b_1 _12339_ (.A_N(net27),
    .B(net26),
    .X(_05107_));
 sky130_fd_sc_hd__a221o_1 _12340_ (.A1(net41),
    .A2(_05084_),
    .B1(_05107_),
    .B2(net43),
    .C1(net29),
    .X(_05108_));
 sky130_fd_sc_hd__o21ai_1 _12341_ (.A1(_05100_),
    .A2(_05106_),
    .B1(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__o22a_1 _12342_ (.A1(_05101_),
    .A2(_05105_),
    .B1(_05109_),
    .B2(net28),
    .X(_05110_));
 sky130_fd_sc_hd__a22oi_1 _12343_ (.A1(_04323_),
    .A2(_05084_),
    .B1(_05107_),
    .B2(net68),
    .Y(_05111_));
 sky130_fd_sc_hd__and4_1 _12344_ (.A(_05082_),
    .B(_05083_),
    .C(_04021_),
    .D(_05085_),
    .X(_05112_));
 sky130_fd_sc_hd__a31o_1 _12345_ (.A1(net42),
    .A2(_05103_),
    .A3(_05085_),
    .B1(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__o21ba_1 _12346_ (.A1(_05101_),
    .A2(_05111_),
    .B1_N(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__a221oi_2 _12347_ (.A1(_05090_),
    .A2(_05102_),
    .B1(_05110_),
    .B2(_05114_),
    .C1(net30),
    .Y(_05115_));
 sky130_fd_sc_hd__mux4_1 _12348_ (.A0(_03473_),
    .A1(_04814_),
    .A2(_04317_),
    .A3(_04809_),
    .S0(_05083_),
    .S1(_05082_),
    .X(_05116_));
 sky130_fd_sc_hd__a31o_1 _12349_ (.A1(net29),
    .A2(net28),
    .A3(_05116_),
    .B1(net30),
    .X(_05117_));
 sky130_fd_sc_hd__mux4_1 _12350_ (.A0(_04813_),
    .A1(_04811_),
    .A2(_04006_),
    .A3(_03475_),
    .S0(_05083_),
    .S1(_05082_),
    .X(_05118_));
 sky130_fd_sc_hd__or2_1 _12351_ (.A(net28),
    .B(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__mux2_1 _12352_ (.A0(_04154_),
    .A1(_03477_),
    .S(_05087_),
    .X(_05120_));
 sky130_fd_sc_hd__o21ai_1 _12353_ (.A1(net29),
    .A2(_05094_),
    .B1(net30),
    .Y(_05121_));
 sky130_fd_sc_hd__o211a_1 _12354_ (.A1(_05101_),
    .A2(_05120_),
    .B1(_05121_),
    .C1(net31),
    .X(_05122_));
 sky130_fd_sc_hd__and3_1 _12355_ (.A(_05117_),
    .B(_05119_),
    .C(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__a2111oi_2 _12356_ (.A1(net124),
    .A2(_05082_),
    .B1(_05087_),
    .C1(net29),
    .D1(net28),
    .Y(_05124_));
 sky130_fd_sc_hd__a22o_1 _12357_ (.A1(net49),
    .A2(_05084_),
    .B1(_05107_),
    .B2(net50),
    .X(_05125_));
 sky130_fd_sc_hd__a21oi_1 _12358_ (.A1(net52),
    .A2(_05103_),
    .B1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__clkinv_2 _12359_ (.A(\gpout4.clk_div[1] ),
    .Y(_05127_));
 sky130_fd_sc_hd__a2bb2o_1 _12360_ (.A1_N(_05127_),
    .A2_N(_05099_),
    .B1(_05107_),
    .B2(net1),
    .X(_05128_));
 sky130_fd_sc_hd__a2bb2o_1 _12361_ (.A1_N(_05101_),
    .A2_N(_05126_),
    .B1(_05128_),
    .B2(_05085_),
    .X(_05129_));
 sky130_fd_sc_hd__o21a_2 _12362_ (.A1(_05124_),
    .A2(_05129_),
    .B1(_05081_),
    .X(_05130_));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(_04883_),
    .A1(_04884_),
    .S(_05083_),
    .X(_05131_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(_04886_),
    .A1(_04887_),
    .S(_05083_),
    .X(_05132_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(_04989_),
    .A1(_04990_),
    .S(_05083_),
    .X(_05133_));
 sky130_fd_sc_hd__mux4_1 _12366_ (.A0(_04891_),
    .A1(_04992_),
    .A2(_04890_),
    .A3(_04892_),
    .S0(_05091_),
    .S1(_05083_),
    .X(_05134_));
 sky130_fd_sc_hd__mux4_1 _12367_ (.A0(_05131_),
    .A1(_05132_),
    .A2(_05133_),
    .A3(_05134_),
    .S0(net28),
    .S1(_05082_),
    .X(_05135_));
 sky130_fd_sc_hd__and3b_1 _12368_ (.A_N(_05121_),
    .B(_05135_),
    .C(net31),
    .X(_05136_));
 sky130_fd_sc_hd__or4_2 _12369_ (.A(_05115_),
    .B(_05123_),
    .C(_05130_),
    .D(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__o2bb2a_2 _12370_ (.A1_N(_04738_),
    .A2_N(_05086_),
    .B1(_05098_),
    .B2(_05137_),
    .X(net57));
 sky130_fd_sc_hd__nor3_2 _12371_ (.A(net35),
    .B(net36),
    .C(net37),
    .Y(_05138_));
 sky130_fd_sc_hd__nor2_2 _12372_ (.A(net33),
    .B(net32),
    .Y(_05139_));
 sky130_fd_sc_hd__nor3b_1 _12373_ (.A(net34),
    .B(net64),
    .C_N(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__inv_2 _12374_ (.A(net33),
    .Y(_05141_));
 sky130_fd_sc_hd__and2_1 _12375_ (.A(_05141_),
    .B(net32),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_4 _12376_ (.A(net32),
    .X(_05143_));
 sky130_fd_sc_hd__nor2_1 _12377_ (.A(_05141_),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__clkbuf_4 _12378_ (.A(net33),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_4 _12379_ (.A(_05143_),
    .X(_05146_));
 sky130_fd_sc_hd__and3_1 _12380_ (.A(_04867_),
    .B(_05145_),
    .C(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__a221o_1 _12381_ (.A1(net52),
    .A2(_05144_),
    .B1(_05139_),
    .B2(net49),
    .C1(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__inv_2 _12382_ (.A(net34),
    .Y(_05149_));
 sky130_fd_sc_hd__a211o_1 _12383_ (.A1(net50),
    .A2(_05142_),
    .B1(_05148_),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a21oi_2 _12384_ (.A1(net123),
    .A2(_05145_),
    .B1(_05146_),
    .Y(_05151_));
 sky130_fd_sc_hd__a311o_2 _12385_ (.A1(_05145_),
    .A2(_05146_),
    .A3(\gpout5.clk_div[1] ),
    .B1(_05151_),
    .C1(net34),
    .X(_05152_));
 sky130_fd_sc_hd__inv_2 _12386_ (.A(net35),
    .Y(_05153_));
 sky130_fd_sc_hd__mux4_1 _12387_ (.A0(_03474_),
    .A1(_04814_),
    .A2(_04317_),
    .A3(_04809_),
    .S0(_05146_),
    .S1(_05145_),
    .X(_05154_));
 sky130_fd_sc_hd__and3_1 _12388_ (.A(net40),
    .B(_05145_),
    .C(_05143_),
    .X(_05155_));
 sky130_fd_sc_hd__a221o_1 _12389_ (.A1(net38),
    .A2(_05142_),
    .B1(_05139_),
    .B2(net48),
    .C1(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__a211o_1 _12390_ (.A1(net39),
    .A2(_05144_),
    .B1(_05156_),
    .C1(_05153_),
    .X(_05157_));
 sky130_fd_sc_hd__a211o_1 _12391_ (.A1(net41),
    .A2(_05139_),
    .B1(net34),
    .C1(net35),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_1 _12392_ (.A1(net43),
    .A2(_05142_),
    .B1(_05144_),
    .B2(net42),
    .C1(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a31o_1 _12393_ (.A1(_05145_),
    .A2(_05143_),
    .A3(_04021_),
    .B1(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__a22o_1 _12394_ (.A1(net46),
    .A2(_05144_),
    .B1(_05139_),
    .B2(_04323_),
    .X(_05161_));
 sky130_fd_sc_hd__a31o_1 _12395_ (.A1(net47),
    .A2(_05145_),
    .A3(_05143_),
    .B1(_05149_),
    .X(_05162_));
 sky130_fd_sc_hd__a211o_1 _12396_ (.A1(net68),
    .A2(_05142_),
    .B1(_05161_),
    .C1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__a32o_1 _12397_ (.A1(_05157_),
    .A2(_05160_),
    .A3(_05163_),
    .B1(net34),
    .B2(net35),
    .X(_05164_));
 sky130_fd_sc_hd__o31a_1 _12398_ (.A1(_05153_),
    .A2(_05149_),
    .A3(_05154_),
    .B1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__mux4_1 _12399_ (.A0(_04006_),
    .A1(_03475_),
    .A2(_04992_),
    .A3(_04892_),
    .S0(_05143_),
    .S1(net34),
    .X(_05166_));
 sky130_fd_sc_hd__mux2_1 _12400_ (.A0(_04154_),
    .A1(_03477_),
    .S(_05143_),
    .X(_05167_));
 sky130_fd_sc_hd__and2_1 _12401_ (.A(net34),
    .B(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(_04813_),
    .A1(_04811_),
    .S(_05143_),
    .X(_05169_));
 sky130_fd_sc_hd__a21o_1 _12403_ (.A1(_05149_),
    .A2(_05169_),
    .B1(_05145_),
    .X(_05170_));
 sky130_fd_sc_hd__o221a_1 _12404_ (.A1(_05141_),
    .A2(_05166_),
    .B1(_05168_),
    .B2(_05170_),
    .C1(_05153_),
    .X(_05171_));
 sky130_fd_sc_hd__mux4_1 _12405_ (.A0(_04989_),
    .A1(\gpout0.vpos[5] ),
    .A2(_04891_),
    .A3(_04890_),
    .S0(_05143_),
    .S1(net34),
    .X(_05172_));
 sky130_fd_sc_hd__mux4_1 _12406_ (.A0(_04883_),
    .A1(_04884_),
    .A2(_04886_),
    .A3(_04887_),
    .S0(_05143_),
    .S1(net34),
    .X(_05173_));
 sky130_fd_sc_hd__or2_1 _12407_ (.A(_05145_),
    .B(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o211a_1 _12408_ (.A1(_05141_),
    .A2(_05172_),
    .B1(_05174_),
    .C1(net35),
    .X(_05175_));
 sky130_fd_sc_hd__or3b_1 _12409_ (.A(_05171_),
    .B(_05175_),
    .C_N(net36),
    .X(_05176_));
 sky130_fd_sc_hd__o211a_1 _12410_ (.A1(net36),
    .A2(_05165_),
    .B1(_05176_),
    .C1(net37),
    .X(_05177_));
 sky130_fd_sc_hd__a31o_2 _12411_ (.A1(_05150_),
    .A2(_05138_),
    .A3(_05152_),
    .B1(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__nand2_1 _12412_ (.A(_05146_),
    .B(_04666_),
    .Y(_05179_));
 sky130_fd_sc_hd__o211a_1 _12413_ (.A1(_05146_),
    .A2(net61),
    .B1(_05179_),
    .C1(net36),
    .X(_05180_));
 sky130_fd_sc_hd__nor2_1 _12414_ (.A(_05146_),
    .B(_04325_),
    .Y(_05181_));
 sky130_fd_sc_hd__a211o_1 _12415_ (.A1(_05146_),
    .A2(net66),
    .B1(_05181_),
    .C1(net36),
    .X(_05182_));
 sky130_fd_sc_hd__nand2_1 _12416_ (.A(_05146_),
    .B(net64),
    .Y(_05183_));
 sky130_fd_sc_hd__o2111a_1 _12417_ (.A1(_05146_),
    .A2(_04738_),
    .B1(_05183_),
    .C1(net35),
    .D1(net36),
    .X(_05184_));
 sky130_fd_sc_hd__and4bb_1 _12418_ (.A_N(net37),
    .B_N(_05184_),
    .C(_05145_),
    .D(net34),
    .X(_05185_));
 sky130_fd_sc_hd__o211a_1 _12419_ (.A1(net35),
    .A2(_05180_),
    .B1(_05182_),
    .C1(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__o2bb2a_2 _12420_ (.A1_N(_05138_),
    .A2_N(_05140_),
    .B1(_05178_),
    .B2(_05186_),
    .X(net58));
 sky130_fd_sc_hd__inv_2 _12421_ (.A(\rbzero.hsync ),
    .Y(net59));
 sky130_fd_sc_hd__and3_1 _12422_ (.A(net71),
    .B(\rbzero.wall_tracer.state[9] ),
    .C(_03480_),
    .X(_05187_));
 sky130_fd_sc_hd__buf_2 _12423_ (.A(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__clkbuf_4 _12424_ (.A(_05188_),
    .X(_00004_));
 sky130_fd_sc_hd__nor2_1 _12425_ (.A(_04032_),
    .B(_03914_),
    .Y(_00005_));
 sky130_fd_sc_hd__buf_4 _12426_ (.A(_03480_),
    .X(_05189_));
 sky130_fd_sc_hd__buf_6 _12427_ (.A(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__and3_1 _12428_ (.A(net71),
    .B(\rbzero.wall_tracer.state[12] ),
    .C(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__clkbuf_1 _12429_ (.A(_05191_),
    .X(_00001_));
 sky130_fd_sc_hd__and3_1 _12430_ (.A(net71),
    .B(\rbzero.wall_tracer.state[7] ),
    .C(_05190_),
    .X(_05192_));
 sky130_fd_sc_hd__clkbuf_1 _12431_ (.A(_05192_),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_1 _12432_ (.A(_04002_),
    .B(_03914_),
    .Y(_00003_));
 sky130_fd_sc_hd__clkinv_4 _12433_ (.A(\rbzero.wall_tracer.state[3] ),
    .Y(_05193_));
 sky130_fd_sc_hd__buf_4 _12434_ (.A(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__nor2_1 _12435_ (.A(_05194_),
    .B(_03914_),
    .Y(_00007_));
 sky130_fd_sc_hd__buf_4 _12436_ (.A(\rbzero.wall_tracer.state[6] ),
    .X(_05195_));
 sky130_fd_sc_hd__clkinv_4 _12437_ (.A(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__buf_4 _12438_ (.A(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__buf_6 _12439_ (.A(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__nor2_1 _12440_ (.A(_05198_),
    .B(_03914_),
    .Y(_00010_));
 sky130_fd_sc_hd__and3_1 _12441_ (.A(net71),
    .B(\rbzero.wall_tracer.state[5] ),
    .C(_05190_),
    .X(_05199_));
 sky130_fd_sc_hd__clkbuf_1 _12442_ (.A(_05199_),
    .X(_00009_));
 sky130_fd_sc_hd__and3_1 _12443_ (.A(net71),
    .B(\rbzero.wall_tracer.state[4] ),
    .C(_03480_),
    .X(_05200_));
 sky130_fd_sc_hd__buf_2 _12444_ (.A(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__clkbuf_4 _12445_ (.A(_05201_),
    .X(_00008_));
 sky130_fd_sc_hd__and3_1 _12446_ (.A(net71),
    .B(\rbzero.wall_tracer.state[2] ),
    .C(_05190_),
    .X(_05202_));
 sky130_fd_sc_hd__clkbuf_1 _12447_ (.A(_05202_),
    .X(_00006_));
 sky130_fd_sc_hd__buf_6 _12448_ (.A(\rbzero.wall_tracer.state[1] ),
    .X(_05203_));
 sky130_fd_sc_hd__buf_8 _12449_ (.A(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__mux2_1 _12450_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_03925_),
    .S(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__buf_4 _12451_ (.A(_05195_),
    .X(_05206_));
 sky130_fd_sc_hd__buf_4 _12452_ (.A(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__buf_4 _12453_ (.A(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__clkbuf_4 _12454_ (.A(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__buf_4 _12455_ (.A(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__buf_6 _12456_ (.A(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__inv_2 _12457_ (.A(\rbzero.wall_tracer.trackDistX[11] ),
    .Y(_05212_));
 sky130_fd_sc_hd__and2_1 _12458_ (.A(_05212_),
    .B(\rbzero.wall_tracer.trackDistY[11] ),
    .X(_05213_));
 sky130_fd_sc_hd__inv_2 _12459_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .Y(_05214_));
 sky130_fd_sc_hd__inv_2 _12460_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .Y(_05215_));
 sky130_fd_sc_hd__a2bb2o_1 _12461_ (.A1_N(_05214_),
    .A2_N(\rbzero.wall_tracer.trackDistX[10] ),
    .B1(\rbzero.wall_tracer.trackDistY[9] ),
    .B2(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__inv_2 _12462_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .Y(_05217_));
 sky130_fd_sc_hd__inv_2 _12463_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .Y(_05218_));
 sky130_fd_sc_hd__a22o_1 _12464_ (.A1(_05217_),
    .A2(\rbzero.wall_tracer.trackDistY[8] ),
    .B1(\rbzero.wall_tracer.trackDistY[7] ),
    .B2(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__inv_2 _12465_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .Y(_05220_));
 sky130_fd_sc_hd__a2bb2o_1 _12466_ (.A1_N(\rbzero.wall_tracer.trackDistY[7] ),
    .A2_N(_05218_),
    .B1(_05220_),
    .B2(\rbzero.wall_tracer.trackDistX[6] ),
    .X(_05221_));
 sky130_fd_sc_hd__inv_2 _12467_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .Y(_05222_));
 sky130_fd_sc_hd__a2bb2o_1 _12468_ (.A1_N(_05220_),
    .A2_N(\rbzero.wall_tracer.trackDistX[6] ),
    .B1(\rbzero.wall_tracer.trackDistY[5] ),
    .B2(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__inv_2 _12469_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .Y(_05224_));
 sky130_fd_sc_hd__o22ai_1 _12470_ (.A1(\rbzero.wall_tracer.trackDistY[5] ),
    .A2(_05222_),
    .B1(_05224_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .Y(_05225_));
 sky130_fd_sc_hd__and2b_1 _12471_ (.A_N(_05223_),
    .B(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__nor2_1 _12472_ (.A(_05221_),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__o22a_1 _12473_ (.A1(\rbzero.wall_tracer.trackDistY[9] ),
    .A2(_05215_),
    .B1(_05217_),
    .B2(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_05228_));
 sky130_fd_sc_hd__o21a_1 _12474_ (.A1(_05219_),
    .A2(_05227_),
    .B1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__nor2_1 _12475_ (.A(_05212_),
    .B(\rbzero.wall_tracer.trackDistY[11] ),
    .Y(_05230_));
 sky130_fd_sc_hd__a21oi_1 _12476_ (.A1(_05214_),
    .A2(\rbzero.wall_tracer.trackDistX[10] ),
    .B1(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21a_1 _12477_ (.A1(_05216_),
    .A2(_05229_),
    .B1(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__or4_1 _12478_ (.A(_05219_),
    .B(_05221_),
    .C(_05223_),
    .D(_05225_),
    .X(_05233_));
 sky130_fd_sc_hd__or4_1 _12479_ (.A(_05233_),
    .B(_05216_),
    .C(_05213_),
    .D(_05230_),
    .X(_05234_));
 sky130_fd_sc_hd__a221o_1 _12480_ (.A1(_05214_),
    .A2(\rbzero.wall_tracer.trackDistX[10] ),
    .B1(_05224_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .C1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__inv_2 _12481_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .Y(_05236_));
 sky130_fd_sc_hd__inv_2 _12482_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .Y(_05237_));
 sky130_fd_sc_hd__inv_2 _12483_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .Y(_05238_));
 sky130_fd_sc_hd__inv_2 _12484_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .Y(_05239_));
 sky130_fd_sc_hd__inv_2 _12485_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .Y(_05240_));
 sky130_fd_sc_hd__inv_2 _12486_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .Y(_05241_));
 sky130_fd_sc_hd__inv_2 _12487_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .Y(_05242_));
 sky130_fd_sc_hd__inv_2 _12488_ (.A(\rbzero.wall_tracer.trackDistX[-12] ),
    .Y(_05243_));
 sky130_fd_sc_hd__o211a_1 _12489_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(_05242_),
    .B1(\rbzero.wall_tracer.trackDistY[-12] ),
    .C1(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__a221o_1 _12490_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(_05241_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .B2(_05242_),
    .C1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__o221a_1 _12491_ (.A1(\rbzero.wall_tracer.trackDistY[-9] ),
    .A2(_05240_),
    .B1(\rbzero.wall_tracer.trackDistY[-10] ),
    .B2(_05241_),
    .C1(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__a221o_1 _12492_ (.A1(_05239_),
    .A2(\rbzero.wall_tracer.trackDistY[-8] ),
    .B1(\rbzero.wall_tracer.trackDistY[-9] ),
    .B2(_05240_),
    .C1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__o221a_1 _12493_ (.A1(\rbzero.wall_tracer.trackDistY[-7] ),
    .A2(_05238_),
    .B1(_05239_),
    .B2(\rbzero.wall_tracer.trackDistY[-8] ),
    .C1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__a221o_1 _12494_ (.A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .A2(_05237_),
    .B1(\rbzero.wall_tracer.trackDistY[-7] ),
    .B2(_05238_),
    .C1(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__o221a_1 _12495_ (.A1(\rbzero.wall_tracer.trackDistY[-5] ),
    .A2(_05236_),
    .B1(\rbzero.wall_tracer.trackDistY[-6] ),
    .B2(_05237_),
    .C1(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__inv_2 _12496_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .Y(_05251_));
 sky130_fd_sc_hd__inv_2 _12497_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .Y(_05252_));
 sky130_fd_sc_hd__o22a_1 _12498_ (.A1(_05251_),
    .A2(\rbzero.wall_tracer.trackDistX[-2] ),
    .B1(_05252_),
    .B2(\rbzero.wall_tracer.trackDistX[-3] ),
    .X(_05253_));
 sky130_fd_sc_hd__inv_2 _12499_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .Y(_05254_));
 sky130_fd_sc_hd__inv_2 _12500_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .Y(_05255_));
 sky130_fd_sc_hd__o22a_1 _12501_ (.A1(_05254_),
    .A2(\rbzero.wall_tracer.trackDistX[2] ),
    .B1(_05255_),
    .B2(\rbzero.wall_tracer.trackDistX[1] ),
    .X(_05256_));
 sky130_fd_sc_hd__inv_2 _12502_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_05257_));
 sky130_fd_sc_hd__inv_2 _12503_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .Y(_05258_));
 sky130_fd_sc_hd__o22a_1 _12504_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(_05257_),
    .B1(_05258_),
    .B2(\rbzero.wall_tracer.trackDistX[-1] ),
    .X(_05259_));
 sky130_fd_sc_hd__nand3_1 _12505_ (.A(_05253_),
    .B(_05256_),
    .C(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__a22o_1 _12506_ (.A1(_05255_),
    .A2(\rbzero.wall_tracer.trackDistX[1] ),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_05257_),
    .X(_05261_));
 sky130_fd_sc_hd__a22o_1 _12507_ (.A1(_05258_),
    .A2(\rbzero.wall_tracer.trackDistX[-1] ),
    .B1(_05251_),
    .B2(\rbzero.wall_tracer.trackDistX[-2] ),
    .X(_05262_));
 sky130_fd_sc_hd__inv_2 _12508_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .Y(_05263_));
 sky130_fd_sc_hd__inv_2 _12509_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .Y(_05264_));
 sky130_fd_sc_hd__a22o_1 _12510_ (.A1(\rbzero.wall_tracer.trackDistY[3] ),
    .A2(_05264_),
    .B1(\rbzero.wall_tracer.trackDistY[-5] ),
    .B2(_05236_),
    .X(_05265_));
 sky130_fd_sc_hd__a21o_1 _12511_ (.A1(_05263_),
    .A2(\rbzero.wall_tracer.trackDistY[-4] ),
    .B1(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__inv_2 _12512_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .Y(_05267_));
 sky130_fd_sc_hd__inv_2 _12513_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .Y(_05268_));
 sky130_fd_sc_hd__o22a_1 _12514_ (.A1(\rbzero.wall_tracer.trackDistY[3] ),
    .A2(_05264_),
    .B1(\rbzero.wall_tracer.trackDistY[2] ),
    .B2(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__o221a_1 _12515_ (.A1(\rbzero.wall_tracer.trackDistY[-3] ),
    .A2(_05267_),
    .B1(_05263_),
    .B2(\rbzero.wall_tracer.trackDistY[-4] ),
    .C1(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__or4b_1 _12516_ (.A(_05261_),
    .B(_05262_),
    .C(_05266_),
    .D_N(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__a2bb2o_1 _12517_ (.A1_N(_05263_),
    .A2_N(\rbzero.wall_tracer.trackDistY[-4] ),
    .B1(_05252_),
    .B2(\rbzero.wall_tracer.trackDistX[-3] ),
    .X(_05272_));
 sky130_fd_sc_hd__a211o_1 _12518_ (.A1(_05272_),
    .A2(_05253_),
    .B1(_05261_),
    .C1(_05262_),
    .X(_05273_));
 sky130_fd_sc_hd__o211ai_1 _12519_ (.A1(_05261_),
    .A2(_05259_),
    .B1(_05256_),
    .C1(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__a22o_1 _12520_ (.A1(\rbzero.wall_tracer.trackDistY[3] ),
    .A2(_05264_),
    .B1(_05269_),
    .B2(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__o31a_1 _12521_ (.A1(_05250_),
    .A2(_05260_),
    .A3(_05271_),
    .B1(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__or3b_1 _12522_ (.A(_05235_),
    .B(_05276_),
    .C_N(_05228_),
    .X(_05277_));
 sky130_fd_sc_hd__o21a_4 _12523_ (.A1(_05213_),
    .A2(_05232_),
    .B1(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__inv_2 _12524_ (.A(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__nor2_1 _12525_ (.A(_03968_),
    .B(_03998_),
    .Y(_05280_));
 sky130_fd_sc_hd__nor2_1 _12526_ (.A(_03912_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__o211a_1 _12527_ (.A1(_04017_),
    .A2(_05279_),
    .B1(_05281_),
    .C1(_03970_),
    .X(_05282_));
 sky130_fd_sc_hd__o21ai_4 _12528_ (.A1(_05203_),
    .A2(_05211_),
    .B1(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__clkbuf_4 _12529_ (.A(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__mux2_1 _12530_ (.A0(_05205_),
    .A1(\rbzero.map_rom.d6 ),
    .S(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_1 _12531_ (.A(_05285_),
    .X(_00401_));
 sky130_fd_sc_hd__or2_1 _12532_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_05286_));
 sky130_fd_sc_hd__and2_1 _12533_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_05287_));
 sky130_fd_sc_hd__a31o_1 _12534_ (.A1(\rbzero.debug_overlay.facingY[-1] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .A3(_05286_),
    .B1(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__or2_2 _12535_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_05289_));
 sky130_fd_sc_hd__or2_1 _12536_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_05290_));
 sky130_fd_sc_hd__xor2_2 _12537_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_05291_));
 sky130_fd_sc_hd__and2_1 _12538_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_05292_));
 sky130_fd_sc_hd__a31o_1 _12539_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_05291_),
    .B1(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__and2_1 _12540_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_05294_));
 sky130_fd_sc_hd__a221o_2 _12541_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_05290_),
    .B2(_05293_),
    .C1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__xor2_1 _12542_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_05296_));
 sky130_fd_sc_hd__nand2_1 _12543_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_05297_));
 sky130_fd_sc_hd__or2_1 _12544_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_05298_));
 sky130_fd_sc_hd__and2_1 _12545_ (.A(_05297_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__and2_1 _12546_ (.A(_05296_),
    .B(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__and2_1 _12547_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_05301_));
 sky130_fd_sc_hd__nor2_1 _12548_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_05302_));
 sky130_fd_sc_hd__nor2_1 _12549_ (.A(_05301_),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nor2_1 _12550_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_05304_));
 sky130_fd_sc_hd__and2_1 _12551_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_05305_));
 sky130_fd_sc_hd__nor2_1 _12552_ (.A(_05304_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__and2_1 _12553_ (.A(_05303_),
    .B(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__and4_1 _12554_ (.A(_05289_),
    .B(_05295_),
    .C(_05300_),
    .D(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__or2_1 _12555_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_05309_));
 sky130_fd_sc_hd__o21a_1 _12556_ (.A1(_05301_),
    .A2(_05305_),
    .B1(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__o211a_1 _12557_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[6] ),
    .B1(\rbzero.wall_tracer.rayAddendY[5] ),
    .C1(\rbzero.debug_overlay.facingY[-3] ),
    .X(_05311_));
 sky130_fd_sc_hd__a221o_1 _12558_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[6] ),
    .B1(_05300_),
    .B2(_05310_),
    .C1(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__nor2_1 _12559_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_05313_));
 sky130_fd_sc_hd__nor2_1 _12560_ (.A(_05313_),
    .B(_05287_),
    .Y(_05314_));
 sky130_fd_sc_hd__and2_1 _12561_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_05315_));
 sky130_fd_sc_hd__nor2_1 _12562_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_05316_));
 sky130_fd_sc_hd__or2_1 _12563_ (.A(_05315_),
    .B(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__inv_2 _12564_ (.A(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__o211a_1 _12565_ (.A1(_05308_),
    .A2(_05312_),
    .B1(_05314_),
    .C1(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__xor2_1 _12566_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_05320_));
 sky130_fd_sc_hd__or2_1 _12567_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_05321_));
 sky130_fd_sc_hd__nand2_1 _12568_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_05322_));
 sky130_fd_sc_hd__and2_1 _12569_ (.A(_05321_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__o211ai_2 _12570_ (.A1(_05288_),
    .A2(_05319_),
    .B1(_05320_),
    .C1(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__o21ai_1 _12571_ (.A1(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2(\rbzero.wall_tracer.rayAddendY[9] ),
    .B1(\rbzero.debug_overlay.facingY[10] ),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _12572_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[11] ),
    .Y(_05326_));
 sky130_fd_sc_hd__or2_1 _12573_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[11] ),
    .X(_05327_));
 sky130_fd_sc_hd__and2_1 _12574_ (.A(_05326_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__a21o_1 _12575_ (.A1(_05324_),
    .A2(_05325_),
    .B1(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__nand3_1 _12576_ (.A(_05324_),
    .B(_05325_),
    .C(_05328_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _12577_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__o21ai_1 _12578_ (.A1(_05288_),
    .A2(_05319_),
    .B1(_05323_),
    .Y(_05332_));
 sky130_fd_sc_hd__and3_1 _12579_ (.A(_05320_),
    .B(_05322_),
    .C(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__a21oi_1 _12580_ (.A1(_05322_),
    .A2(_05332_),
    .B1(_05320_),
    .Y(_05334_));
 sky130_fd_sc_hd__or2_1 _12581_ (.A(_05333_),
    .B(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__and3_1 _12582_ (.A(_05289_),
    .B(_05295_),
    .C(_05303_),
    .X(_05336_));
 sky130_fd_sc_hd__o311ai_4 _12583_ (.A1(_05301_),
    .A2(_05336_),
    .A3(_05305_),
    .B1(_05309_),
    .C1(_05299_),
    .Y(_05337_));
 sky130_fd_sc_hd__a21bo_1 _12584_ (.A1(_05297_),
    .A2(_05337_),
    .B1_N(_05296_),
    .X(_05338_));
 sky130_fd_sc_hd__nand3b_1 _12585_ (.A_N(_05296_),
    .B(_05297_),
    .C(_05337_),
    .Y(_05339_));
 sky130_fd_sc_hd__and2_1 _12586_ (.A(_05338_),
    .B(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__or3_1 _12587_ (.A(_05323_),
    .B(_05288_),
    .C(_05319_),
    .X(_05341_));
 sky130_fd_sc_hd__and2_1 _12588_ (.A(_05332_),
    .B(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__a31o_1 _12589_ (.A1(_05289_),
    .A2(_05295_),
    .A3(_05303_),
    .B1(_05301_),
    .X(_05343_));
 sky130_fd_sc_hd__a211o_1 _12590_ (.A1(_05309_),
    .A2(_05343_),
    .B1(_05305_),
    .C1(_05299_),
    .X(_05344_));
 sky130_fd_sc_hd__and2_1 _12591_ (.A(_05337_),
    .B(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__xor2_1 _12592_ (.A(_05306_),
    .B(_05343_),
    .X(_05346_));
 sky130_fd_sc_hd__nand3_1 _12593_ (.A(_05289_),
    .B(_05295_),
    .C(_05303_),
    .Y(_05347_));
 sky130_fd_sc_hd__a21o_1 _12594_ (.A1(_05289_),
    .A2(_05295_),
    .B1(_05303_),
    .X(_05348_));
 sky130_fd_sc_hd__and2_1 _12595_ (.A(_05347_),
    .B(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__and2b_1 _12596_ (.A_N(_05294_),
    .B(_05290_),
    .X(_05350_));
 sky130_fd_sc_hd__xor2_1 _12597_ (.A(_05350_),
    .B(_05293_),
    .X(_05351_));
 sky130_fd_sc_hd__nand2_1 _12598_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_05352_));
 sky130_fd_sc_hd__xnor2_2 _12599_ (.A(_05352_),
    .B(_05291_),
    .Y(_05353_));
 sky130_fd_sc_hd__or2_1 _12600_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_05354_));
 sky130_fd_sc_hd__and2_1 _12601_ (.A(_05352_),
    .B(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__or4_1 _12602_ (.A(\rbzero.wall_tracer.rayAddendY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .C(\rbzero.wall_tracer.rayAddendY[-2] ),
    .D(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__nand2_1 _12603_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_05357_));
 sky130_fd_sc_hd__nand2_1 _12604_ (.A(_05289_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__a21o_1 _12605_ (.A1(_05290_),
    .A2(_05293_),
    .B1(_05294_),
    .X(_05359_));
 sky130_fd_sc_hd__xnor2_2 _12606_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__or4_1 _12607_ (.A(_05351_),
    .B(_05353_),
    .C(_05356_),
    .D(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__o21ai_1 _12608_ (.A1(_05308_),
    .A2(_05312_),
    .B1(_05318_),
    .Y(_05362_));
 sky130_fd_sc_hd__or3_1 _12609_ (.A(_05318_),
    .B(_05308_),
    .C(_05312_),
    .X(_05363_));
 sky130_fd_sc_hd__and2_1 _12610_ (.A(_05362_),
    .B(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__or4_1 _12611_ (.A(_05346_),
    .B(_05349_),
    .C(_05361_),
    .D(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__o21a_1 _12612_ (.A1(_05308_),
    .A2(_05312_),
    .B1(_05318_),
    .X(_05366_));
 sky130_fd_sc_hd__o21ai_1 _12613_ (.A1(_05315_),
    .A2(_05366_),
    .B1(_05314_),
    .Y(_05367_));
 sky130_fd_sc_hd__or3_1 _12614_ (.A(_05315_),
    .B(_05366_),
    .C(_05314_),
    .X(_05368_));
 sky130_fd_sc_hd__nand2_1 _12615_ (.A(_05367_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__or4b_2 _12616_ (.A(_05342_),
    .B(_05345_),
    .C(_05365_),
    .D_N(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__a21bo_1 _12617_ (.A1(_05324_),
    .A2(_05325_),
    .B1_N(_05326_),
    .X(_05371_));
 sky130_fd_sc_hd__nand2_2 _12618_ (.A(_05327_),
    .B(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__o41ai_4 _12619_ (.A1(_05331_),
    .A2(_05335_),
    .A3(_05340_),
    .A4(_05370_),
    .B1(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__clkbuf_4 _12620_ (.A(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__and2_1 _12621_ (.A(\rbzero.map_rom.c6 ),
    .B(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__nor2_1 _12622_ (.A(_03942_),
    .B(_05374_),
    .Y(_05376_));
 sky130_fd_sc_hd__nor2_1 _12623_ (.A(_05375_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__xnor2_1 _12624_ (.A(_03925_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(\rbzero.debug_overlay.playerY[1] ),
    .A1(_05378_),
    .S(_05204_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _12626_ (.A0(_05379_),
    .A1(_03942_),
    .S(_05284_),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_1 _12627_ (.A(_05380_),
    .X(_00402_));
 sky130_fd_sc_hd__and2_1 _12628_ (.A(\rbzero.map_rom.b6 ),
    .B(_05374_),
    .X(_05381_));
 sky130_fd_sc_hd__nor2_1 _12629_ (.A(_03933_),
    .B(_05374_),
    .Y(_05382_));
 sky130_fd_sc_hd__nor2_1 _12630_ (.A(_05381_),
    .B(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__a21oi_1 _12631_ (.A1(\rbzero.map_rom.d6 ),
    .A2(_05377_),
    .B1(_05375_),
    .Y(_05384_));
 sky130_fd_sc_hd__xnor2_1 _12632_ (.A(_05383_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__mux2_1 _12633_ (.A0(\rbzero.debug_overlay.playerY[2] ),
    .A1(_05385_),
    .S(_05204_),
    .X(_05386_));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(_05386_),
    .A1(_03933_),
    .S(_05284_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _12635_ (.A(_05387_),
    .X(_00403_));
 sky130_fd_sc_hd__or2_1 _12636_ (.A(\rbzero.map_rom.a6 ),
    .B(_05374_),
    .X(_05388_));
 sky130_fd_sc_hd__and2_1 _12637_ (.A(\rbzero.map_rom.a6 ),
    .B(_05374_),
    .X(_05389_));
 sky130_fd_sc_hd__inv_2 _12638_ (.A(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(_05388_),
    .B(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__o21bai_1 _12640_ (.A1(_05382_),
    .A2(_05384_),
    .B1_N(_05381_),
    .Y(_05392_));
 sky130_fd_sc_hd__xnor2_1 _12641_ (.A(_05391_),
    .B(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__buf_4 _12642_ (.A(_05203_),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _12643_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_05393_),
    .S(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__mux2_1 _12644_ (.A0(_05395_),
    .A1(\rbzero.map_rom.a6 ),
    .S(_05284_),
    .X(_05396_));
 sky130_fd_sc_hd__clkbuf_1 _12645_ (.A(_05396_),
    .X(_00404_));
 sky130_fd_sc_hd__clkbuf_4 _12646_ (.A(_05374_),
    .X(_05397_));
 sky130_fd_sc_hd__xnor2_1 _12647_ (.A(_03935_),
    .B(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__or2_1 _12648_ (.A(_05389_),
    .B(_05392_),
    .X(_05399_));
 sky130_fd_sc_hd__nand2_1 _12649_ (.A(_05388_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__xnor2_1 _12650_ (.A(_05398_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__mux2_1 _12651_ (.A0(\rbzero.debug_overlay.playerY[4] ),
    .A1(_05401_),
    .S(_05394_),
    .X(_05402_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(_05402_),
    .A1(\rbzero.map_rom.i_row[4] ),
    .S(_05283_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _12653_ (.A(_05403_),
    .X(_00405_));
 sky130_fd_sc_hd__clkbuf_4 _12654_ (.A(_05397_),
    .X(_05404_));
 sky130_fd_sc_hd__xnor2_1 _12655_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__a32o_1 _12656_ (.A1(_05388_),
    .A2(_05398_),
    .A3(_05399_),
    .B1(_05397_),
    .B2(\rbzero.map_rom.i_row[4] ),
    .X(_05406_));
 sky130_fd_sc_hd__xnor2_1 _12657_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(\rbzero.debug_overlay.playerY[5] ),
    .A1(_05407_),
    .S(_05394_),
    .X(_05408_));
 sky130_fd_sc_hd__mux2_1 _12659_ (.A0(_05408_),
    .A1(\rbzero.wall_tracer.mapY[5] ),
    .S(_05283_),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _12660_ (.A(_05409_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_03919_),
    .S(_05394_),
    .X(_05410_));
 sky130_fd_sc_hd__inv_2 _12662_ (.A(_03999_),
    .Y(_05411_));
 sky130_fd_sc_hd__o221ai_4 _12663_ (.A1(\rbzero.wall_tracer.state[1] ),
    .A2(_05211_),
    .B1(_04017_),
    .B2(_05278_),
    .C1(_05281_),
    .Y(_05412_));
 sky130_fd_sc_hd__nor2_8 _12664_ (.A(_05411_),
    .B(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__buf_6 _12665_ (.A(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__mux2_1 _12666_ (.A0(\rbzero.map_rom.f4 ),
    .A1(_05410_),
    .S(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__clkbuf_1 _12667_ (.A(_05415_),
    .X(_00407_));
 sky130_fd_sc_hd__nand2_1 _12668_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_05416_));
 sky130_fd_sc_hd__or2_1 _12669_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_05417_));
 sky130_fd_sc_hd__nand2_1 _12670_ (.A(_05416_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__nor2_1 _12671_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_1 _12672_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_05420_));
 sky130_fd_sc_hd__and2b_1 _12673_ (.A_N(_05419_),
    .B(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__nor2_1 _12674_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_05422_));
 sky130_fd_sc_hd__nor2_1 _12675_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_05423_));
 sky130_fd_sc_hd__nand2_2 _12676_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_05424_));
 sky130_fd_sc_hd__nor2_1 _12677_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _12678_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _12679_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_05427_));
 sky130_fd_sc_hd__o211a_1 _12680_ (.A1(_05424_),
    .A2(_05425_),
    .B1(_05426_),
    .C1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _12681_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_05429_));
 sky130_fd_sc_hd__o31ai_4 _12682_ (.A1(_05422_),
    .A2(_05423_),
    .A3(_05428_),
    .B1(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _12683_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_05431_));
 sky130_fd_sc_hd__or2_1 _12684_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_05432_));
 sky130_fd_sc_hd__and2_1 _12685_ (.A(_05431_),
    .B(_05432_),
    .X(_05433_));
 sky130_fd_sc_hd__or2_1 _12686_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_05434_));
 sky130_fd_sc_hd__and3_1 _12687_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .C(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__and2_1 _12688_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_05436_));
 sky130_fd_sc_hd__a21o_1 _12689_ (.A1(_05420_),
    .A2(_05431_),
    .B1(_05419_),
    .X(_05437_));
 sky130_fd_sc_hd__or3b_1 _12690_ (.A(_05435_),
    .B(_05436_),
    .C_N(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__a31o_1 _12691_ (.A1(_05421_),
    .A2(_05430_),
    .A3(_05433_),
    .B1(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__or2_1 _12692_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_05440_));
 sky130_fd_sc_hd__o21a_1 _12693_ (.A1(_05436_),
    .A2(_05440_),
    .B1(_05434_),
    .X(_05441_));
 sky130_fd_sc_hd__nand3b_1 _12694_ (.A_N(_05418_),
    .B(_05439_),
    .C(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_1 _12695_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_05443_));
 sky130_fd_sc_hd__nor2_1 _12696_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_05444_));
 sky130_fd_sc_hd__xnor2_2 _12697_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_05445_));
 sky130_fd_sc_hd__a311o_1 _12698_ (.A1(_05416_),
    .A2(_05442_),
    .A3(_05443_),
    .B1(_05444_),
    .C1(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__xnor2_4 _12699_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_05447_));
 sky130_fd_sc_hd__or2_1 _12700_ (.A(\rbzero.wall_tracer.rayAddendX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_05448_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__o21a_1 _12702_ (.A1(_05446_),
    .A2(_05447_),
    .B1(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__or2_1 _12703_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[11] ),
    .X(_05451_));
 sky130_fd_sc_hd__nand2_1 _12704_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[11] ),
    .Y(_05452_));
 sky130_fd_sc_hd__nand2_1 _12705_ (.A(_05451_),
    .B(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__xnor2_2 _12706_ (.A(_05450_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__a21bo_1 _12707_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(\rbzero.wall_tracer.rayAddendX[9] ),
    .B1_N(_05446_),
    .X(_05455_));
 sky130_fd_sc_hd__xor2_4 _12708_ (.A(_05447_),
    .B(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__or2b_1 _12709_ (.A(_05444_),
    .B_N(_05443_),
    .X(_05457_));
 sky130_fd_sc_hd__nand2_1 _12710_ (.A(_05416_),
    .B(_05442_),
    .Y(_05458_));
 sky130_fd_sc_hd__xnor2_2 _12711_ (.A(_05457_),
    .B(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__a21bo_1 _12712_ (.A1(_05439_),
    .A2(_05441_),
    .B1_N(_05418_),
    .X(_05460_));
 sky130_fd_sc_hd__and2_1 _12713_ (.A(_05442_),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__nand2_1 _12714_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_05462_));
 sky130_fd_sc_hd__nand2_1 _12715_ (.A(_05462_),
    .B(_05440_),
    .Y(_05463_));
 sky130_fd_sc_hd__inv_2 _12716_ (.A(_05437_),
    .Y(_05464_));
 sky130_fd_sc_hd__a31o_1 _12717_ (.A1(_05421_),
    .A2(_05430_),
    .A3(_05433_),
    .B1(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__xnor2_2 _12718_ (.A(_05463_),
    .B(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21boi_1 _12719_ (.A1(_05430_),
    .A2(_05433_),
    .B1_N(_05431_),
    .Y(_05467_));
 sky130_fd_sc_hd__xnor2_1 _12720_ (.A(_05421_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__xor2_2 _12721_ (.A(_05430_),
    .B(_05433_),
    .X(_05469_));
 sky130_fd_sc_hd__or2_1 _12722_ (.A(_05423_),
    .B(_05428_),
    .X(_05470_));
 sky130_fd_sc_hd__and2b_1 _12723_ (.A_N(_05422_),
    .B(_05429_),
    .X(_05471_));
 sky130_fd_sc_hd__xnor2_2 _12724_ (.A(_05470_),
    .B(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__o21a_1 _12725_ (.A1(_05424_),
    .A2(_05425_),
    .B1(_05427_),
    .X(_05473_));
 sky130_fd_sc_hd__and2b_1 _12726_ (.A_N(_05423_),
    .B(_05426_),
    .X(_05474_));
 sky130_fd_sc_hd__xnor2_2 _12727_ (.A(_05473_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__or2_1 _12728_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_05476_));
 sky130_fd_sc_hd__and2_1 _12729_ (.A(_05424_),
    .B(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__or4_1 _12730_ (.A(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .C(\rbzero.wall_tracer.rayAddendX[-2] ),
    .D(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__and2_1 _12731_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_05479_));
 sky130_fd_sc_hd__nor2_2 _12732_ (.A(_05479_),
    .B(_05425_),
    .Y(_05480_));
 sky130_fd_sc_hd__xnor2_4 _12733_ (.A(_05424_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__or4_1 _12734_ (.A(_05472_),
    .B(_05475_),
    .C(_05478_),
    .D(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__or4_1 _12735_ (.A(_05466_),
    .B(_05468_),
    .C(_05469_),
    .D(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__nor2_1 _12736_ (.A(_05461_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__nand2_1 _12737_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2_1 _12738_ (.A(_05434_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__a21boi_1 _12739_ (.A1(_05440_),
    .A2(_05465_),
    .B1_N(_05462_),
    .Y(_05487_));
 sky130_fd_sc_hd__xnor2_2 _12740_ (.A(_05486_),
    .B(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__a31o_1 _12741_ (.A1(_05416_),
    .A2(_05442_),
    .A3(_05443_),
    .B1(_05444_),
    .X(_05489_));
 sky130_fd_sc_hd__xnor2_2 _12742_ (.A(_05445_),
    .B(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__and4b_1 _12743_ (.A_N(_05459_),
    .B(_05484_),
    .C(_05488_),
    .D(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__and2_1 _12744_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[11] ),
    .X(_05492_));
 sky130_fd_sc_hd__o211a_1 _12745_ (.A1(_05446_),
    .A2(_05447_),
    .B1(_05451_),
    .C1(_05449_),
    .X(_05493_));
 sky130_fd_sc_hd__or2_2 _12746_ (.A(_05492_),
    .B(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__a31o_4 _12747_ (.A1(_05454_),
    .A2(_05456_),
    .A3(_05491_),
    .B1(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__buf_4 _12748_ (.A(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__xnor2_1 _12749_ (.A(_03924_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__or2_1 _12750_ (.A(\rbzero.map_rom.f4 ),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__nand2_1 _12751_ (.A(\rbzero.map_rom.f4 ),
    .B(_05497_),
    .Y(_05499_));
 sky130_fd_sc_hd__nor2_1 _12752_ (.A(_03926_),
    .B(_05394_),
    .Y(_05500_));
 sky130_fd_sc_hd__a31o_1 _12753_ (.A1(_05204_),
    .A2(_05498_),
    .A3(_05499_),
    .B1(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _12754_ (.A0(\rbzero.map_rom.f3 ),
    .A1(_05501_),
    .S(_05414_),
    .X(_05502_));
 sky130_fd_sc_hd__clkbuf_1 _12755_ (.A(_05502_),
    .X(_00408_));
 sky130_fd_sc_hd__inv_2 _12756_ (.A(_05496_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor2_1 _12757_ (.A(_03929_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__nor2_1 _12758_ (.A(\rbzero.map_rom.f2 ),
    .B(_05496_),
    .Y(_05505_));
 sky130_fd_sc_hd__nor2_1 _12759_ (.A(_05504_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_1 _12760_ (.A1(_03924_),
    .A2(_05503_),
    .B1(_05499_),
    .Y(_05507_));
 sky130_fd_sc_hd__xor2_1 _12761_ (.A(_05506_),
    .B(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(\rbzero.debug_overlay.playerX[2] ),
    .A1(_05508_),
    .S(_05394_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _12763_ (.A0(\rbzero.map_rom.f2 ),
    .A1(_05509_),
    .S(_05414_),
    .X(_05510_));
 sky130_fd_sc_hd__clkbuf_1 _12764_ (.A(_05510_),
    .X(_00409_));
 sky130_fd_sc_hd__nor2_1 _12765_ (.A(_03936_),
    .B(_05503_),
    .Y(_05511_));
 sky130_fd_sc_hd__buf_2 _12766_ (.A(_05496_),
    .X(_05512_));
 sky130_fd_sc_hd__or2_1 _12767_ (.A(\rbzero.map_rom.f1 ),
    .B(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__or2b_1 _12768_ (.A(_05511_),
    .B_N(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__a21o_1 _12769_ (.A1(_05506_),
    .A2(_05507_),
    .B1(_05504_),
    .X(_05515_));
 sky130_fd_sc_hd__xnor2_1 _12770_ (.A(_05514_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__mux2_1 _12771_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_05516_),
    .S(_05394_),
    .X(_05517_));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(\rbzero.map_rom.f1 ),
    .A1(_05517_),
    .S(_05414_),
    .X(_05518_));
 sky130_fd_sc_hd__clkbuf_1 _12773_ (.A(_05518_),
    .X(_00410_));
 sky130_fd_sc_hd__xor2_1 _12774_ (.A(\rbzero.map_rom.i_col[4] ),
    .B(_05512_),
    .X(_05519_));
 sky130_fd_sc_hd__or2_1 _12775_ (.A(_05511_),
    .B(_05515_),
    .X(_05520_));
 sky130_fd_sc_hd__nand2_1 _12776_ (.A(_05513_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__xnor2_1 _12777_ (.A(_05519_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(\rbzero.debug_overlay.playerX[4] ),
    .A1(_05522_),
    .S(_05394_),
    .X(_05523_));
 sky130_fd_sc_hd__mux2_1 _12779_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_05523_),
    .S(_05414_),
    .X(_05524_));
 sky130_fd_sc_hd__clkbuf_1 _12780_ (.A(_05524_),
    .X(_00411_));
 sky130_fd_sc_hd__clkbuf_4 _12781_ (.A(_05512_),
    .X(_05525_));
 sky130_fd_sc_hd__xnor2_1 _12782_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__a32o_1 _12783_ (.A1(_05513_),
    .A2(_05519_),
    .A3(_05520_),
    .B1(_05512_),
    .B2(\rbzero.map_rom.i_col[4] ),
    .X(_05527_));
 sky130_fd_sc_hd__xnor2_1 _12784_ (.A(_05526_),
    .B(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(\rbzero.debug_overlay.playerX[5] ),
    .A1(_05528_),
    .S(_05394_),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _12786_ (.A0(\rbzero.wall_tracer.mapX[5] ),
    .A1(_05529_),
    .S(_05414_),
    .X(_05530_));
 sky130_fd_sc_hd__clkbuf_1 _12787_ (.A(_05530_),
    .X(_00412_));
 sky130_fd_sc_hd__buf_4 _12788_ (.A(_04016_),
    .X(_05531_));
 sky130_fd_sc_hd__buf_6 _12789_ (.A(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__nor2_4 _12790_ (.A(_05532_),
    .B(_05283_),
    .Y(_05533_));
 sky130_fd_sc_hd__xor2_1 _12791_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_05397_),
    .X(_05534_));
 sky130_fd_sc_hd__a21o_1 _12792_ (.A1(\rbzero.wall_tracer.mapY[5] ),
    .A2(_05397_),
    .B1(_05406_),
    .X(_05535_));
 sky130_fd_sc_hd__o21a_1 _12793_ (.A1(\rbzero.wall_tracer.mapY[5] ),
    .A2(_05397_),
    .B1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__or2_1 _12794_ (.A(_05534_),
    .B(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__nand2_1 _12795_ (.A(_05534_),
    .B(_05536_),
    .Y(_05538_));
 sky130_fd_sc_hd__a32o_1 _12796_ (.A1(_05533_),
    .A2(_05537_),
    .A3(_05538_),
    .B1(_05284_),
    .B2(\rbzero.wall_tracer.mapY[6] ),
    .X(_00413_));
 sky130_fd_sc_hd__and2_1 _12797_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_05397_),
    .X(_05539_));
 sky130_fd_sc_hd__a21bo_1 _12798_ (.A1(\rbzero.wall_tracer.mapY[6] ),
    .A2(_05397_),
    .B1_N(_05538_),
    .X(_05540_));
 sky130_fd_sc_hd__o21a_1 _12799_ (.A1(\rbzero.wall_tracer.mapY[7] ),
    .A2(_05397_),
    .B1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__or2b_1 _12800_ (.A(_05539_),
    .B_N(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__nor2_1 _12801_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_05404_),
    .Y(_05543_));
 sky130_fd_sc_hd__o21bai_1 _12802_ (.A1(_05539_),
    .A2(_05543_),
    .B1_N(_05540_),
    .Y(_05544_));
 sky130_fd_sc_hd__a32o_1 _12803_ (.A1(_05533_),
    .A2(_05542_),
    .A3(_05544_),
    .B1(_05284_),
    .B2(\rbzero.wall_tracer.mapY[7] ),
    .X(_00414_));
 sky130_fd_sc_hd__xor2_1 _12804_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_05404_),
    .X(_05545_));
 sky130_fd_sc_hd__or3_1 _12805_ (.A(_05539_),
    .B(_05541_),
    .C(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__o21ai_1 _12806_ (.A1(_05539_),
    .A2(_05541_),
    .B1(_05545_),
    .Y(_05547_));
 sky130_fd_sc_hd__a32o_1 _12807_ (.A1(_05533_),
    .A2(_05546_),
    .A3(_05547_),
    .B1(_05284_),
    .B2(\rbzero.wall_tracer.mapY[8] ),
    .X(_00415_));
 sky130_fd_sc_hd__and2_1 _12808_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_05404_),
    .X(_05548_));
 sky130_fd_sc_hd__nor2_1 _12809_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_05404_),
    .Y(_05549_));
 sky130_fd_sc_hd__a21bo_1 _12810_ (.A1(\rbzero.wall_tracer.mapY[8] ),
    .A2(_05404_),
    .B1_N(_05547_),
    .X(_05550_));
 sky130_fd_sc_hd__o21bai_1 _12811_ (.A1(_05548_),
    .A2(_05549_),
    .B1_N(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__o21a_1 _12812_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_05404_),
    .B1(_05550_),
    .X(_05552_));
 sky130_fd_sc_hd__or2b_1 _12813_ (.A(_05548_),
    .B_N(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__a32o_1 _12814_ (.A1(_05533_),
    .A2(_05551_),
    .A3(_05553_),
    .B1(_05284_),
    .B2(\rbzero.wall_tracer.mapY[9] ),
    .X(_00416_));
 sky130_fd_sc_hd__xor2_1 _12815_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_05404_),
    .X(_05554_));
 sky130_fd_sc_hd__o21ai_1 _12816_ (.A1(_05548_),
    .A2(_05552_),
    .B1(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__or3_1 _12817_ (.A(_05548_),
    .B(_05552_),
    .C(_05554_),
    .X(_05556_));
 sky130_fd_sc_hd__a32o_1 _12818_ (.A1(_05533_),
    .A2(_05555_),
    .A3(_05556_),
    .B1(_05284_),
    .B2(\rbzero.wall_tracer.mapY[10] ),
    .X(_00417_));
 sky130_fd_sc_hd__a21bo_1 _12819_ (.A1(\rbzero.wall_tracer.mapY[10] ),
    .A2(_05404_),
    .B1_N(_05555_),
    .X(_05557_));
 sky130_fd_sc_hd__xnor2_1 _12820_ (.A(\rbzero.wall_tracer.mapY[11] ),
    .B(_05404_),
    .Y(_05558_));
 sky130_fd_sc_hd__xnor2_1 _12821_ (.A(_05557_),
    .B(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__a22o_1 _12822_ (.A1(\rbzero.wall_tracer.mapY[11] ),
    .A2(_05284_),
    .B1(_05533_),
    .B2(_05559_),
    .X(_00418_));
 sky130_fd_sc_hd__clkinv_2 _12823_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_05560_));
 sky130_fd_sc_hd__clkbuf_4 _12824_ (.A(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__or3_2 _12825_ (.A(_05561_),
    .B(_05492_),
    .C(_05493_),
    .X(_05562_));
 sky130_fd_sc_hd__buf_2 _12826_ (.A(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__nor2_1 _12827_ (.A(_03953_),
    .B(_04030_),
    .Y(_05564_));
 sky130_fd_sc_hd__a311o_1 _12828_ (.A1(_04030_),
    .A2(_05327_),
    .A3(_05371_),
    .B1(_05564_),
    .C1(_04001_),
    .X(_05565_));
 sky130_fd_sc_hd__buf_2 _12829_ (.A(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__nand2_2 _12830_ (.A(_05563_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__nor2_1 _12831_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_04031_),
    .Y(_05568_));
 sky130_fd_sc_hd__a211o_1 _12832_ (.A1(_04031_),
    .A2(_05372_),
    .B1(_05568_),
    .C1(_04001_),
    .X(_05569_));
 sky130_fd_sc_hd__inv_2 _12833_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .Y(_05570_));
 sky130_fd_sc_hd__buf_2 _12834_ (.A(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__a31o_1 _12835_ (.A1(_04031_),
    .A2(_05327_),
    .A3(_05371_),
    .B1(_04001_),
    .X(_05572_));
 sky130_fd_sc_hd__a21o_1 _12836_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(_05571_),
    .B1(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__nand2_1 _12837_ (.A(_05563_),
    .B(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__and2_1 _12838_ (.A(_05569_),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__a21o_1 _12839_ (.A1(\rbzero.wall_tracer.visualWallDist[10] ),
    .A2(_05571_),
    .B1(_05572_),
    .X(_05576_));
 sky130_fd_sc_hd__or2_1 _12840_ (.A(_05561_),
    .B(_05468_),
    .X(_05577_));
 sky130_fd_sc_hd__a21o_1 _12841_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_05570_),
    .B1(_04000_),
    .X(_05578_));
 sky130_fd_sc_hd__a21o_1 _12842_ (.A1(_04030_),
    .A2(_05346_),
    .B1(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__and3_1 _12843_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .B(_05347_),
    .C(_05348_),
    .X(_05580_));
 sky130_fd_sc_hd__a21o_1 _12844_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_05570_),
    .B1(_04000_),
    .X(_05581_));
 sky130_fd_sc_hd__o22a_2 _12845_ (.A1(_05561_),
    .A2(_05469_),
    .B1(_05580_),
    .B2(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A1(_05351_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05583_));
 sky130_fd_sc_hd__mux2_2 _12847_ (.A0(_05475_),
    .A1(_05583_),
    .S(_05561_),
    .X(_05584_));
 sky130_fd_sc_hd__or2_1 _12848_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05585_));
 sky130_fd_sc_hd__o211a_1 _12849_ (.A1(_05570_),
    .A2(_05360_),
    .B1(_05585_),
    .C1(_05561_),
    .X(_05586_));
 sky130_fd_sc_hd__and2_1 _12850_ (.A(_04000_),
    .B(_05472_),
    .X(_05587_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05588_));
 sky130_fd_sc_hd__mux2_2 _12852_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_05588_),
    .S(_05560_),
    .X(_05589_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(\rbzero.wall_tracer.visualWallDist[-12] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05590_));
 sky130_fd_sc_hd__mux2_2 _12854_ (.A0(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A1(_05590_),
    .S(_05560_),
    .X(_05591_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05592_));
 sky130_fd_sc_hd__mux2_2 _12856_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_05592_),
    .S(_05560_),
    .X(_05593_));
 sky130_fd_sc_hd__or3_1 _12857_ (.A(_05589_),
    .B(_05591_),
    .C(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_05355_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05595_));
 sky130_fd_sc_hd__mux2_4 _12859_ (.A0(_05477_),
    .A1(_05595_),
    .S(_05560_),
    .X(_05596_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_05353_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_05597_));
 sky130_fd_sc_hd__mux2_2 _12861_ (.A0(_05481_),
    .A1(_05597_),
    .S(_05561_),
    .X(_05598_));
 sky130_fd_sc_hd__nor3_1 _12862_ (.A(_05594_),
    .B(_05596_),
    .C(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__or4b_1 _12863_ (.A(_05584_),
    .B(_05586_),
    .C(_05587_),
    .D_N(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__a211o_2 _12864_ (.A1(_05577_),
    .A2(_05579_),
    .B1(_05582_),
    .C1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__nor2_1 _12865_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_04031_),
    .Y(_05602_));
 sky130_fd_sc_hd__a211o_1 _12866_ (.A1(_04031_),
    .A2(_05372_),
    .B1(_05602_),
    .C1(_04001_),
    .X(_05603_));
 sky130_fd_sc_hd__a21o_1 _12867_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_05571_),
    .B1(_05572_),
    .X(_05604_));
 sky130_fd_sc_hd__nand2_1 _12868_ (.A(_05563_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _12869_ (.A(_05603_),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__a21o_1 _12870_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_05571_),
    .B1(_04000_),
    .X(_05607_));
 sky130_fd_sc_hd__a31o_1 _12871_ (.A1(_04030_),
    .A2(_05367_),
    .A3(_05368_),
    .B1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__o21a_2 _12872_ (.A1(_05561_),
    .A2(_05459_),
    .B1(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__nand2_1 _12873_ (.A(_04000_),
    .B(_05488_),
    .Y(_05610_));
 sky130_fd_sc_hd__a21o_1 _12874_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_05571_),
    .B1(_04000_),
    .X(_05611_));
 sky130_fd_sc_hd__a31o_1 _12875_ (.A1(_04030_),
    .A2(_05338_),
    .A3(_05339_),
    .B1(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__a21o_1 _12876_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_05571_),
    .B1(_04000_),
    .X(_05613_));
 sky130_fd_sc_hd__a31o_1 _12877_ (.A1(_04030_),
    .A2(_05337_),
    .A3(_05344_),
    .B1(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__o21a_2 _12878_ (.A1(_05561_),
    .A2(_05466_),
    .B1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__and3_1 _12879_ (.A(_04030_),
    .B(_05362_),
    .C(_05363_),
    .X(_05616_));
 sky130_fd_sc_hd__a21o_1 _12880_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_05571_),
    .B1(_04000_),
    .X(_05617_));
 sky130_fd_sc_hd__o22a_1 _12881_ (.A1(_05561_),
    .A2(_05461_),
    .B1(_05616_),
    .B2(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__a2111o_1 _12882_ (.A1(_05610_),
    .A2(_05612_),
    .B1(_05615_),
    .C1(_05601_),
    .D1(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__and3_1 _12883_ (.A(_04030_),
    .B(_05332_),
    .C(_05341_),
    .X(_05620_));
 sky130_fd_sc_hd__a21o_1 _12884_ (.A1(\rbzero.wall_tracer.visualWallDist[1] ),
    .A2(_05571_),
    .B1(_04000_),
    .X(_05621_));
 sky130_fd_sc_hd__o2bb2a_2 _12885_ (.A1_N(_04001_),
    .A2_N(_05490_),
    .B1(_05620_),
    .B2(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__or3_1 _12886_ (.A(_05609_),
    .B(_05619_),
    .C(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__o21ai_1 _12887_ (.A1(_05333_),
    .A2(_05334_),
    .B1(_04031_),
    .Y(_05624_));
 sky130_fd_sc_hd__a21oi_1 _12888_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_05571_),
    .B1(_04001_),
    .Y(_05625_));
 sky130_fd_sc_hd__a22oi_4 _12889_ (.A1(_04001_),
    .A2(_05456_),
    .B1(_05624_),
    .B2(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__and2_1 _12890_ (.A(_05562_),
    .B(_05565_),
    .X(_05627_));
 sky130_fd_sc_hd__buf_2 _12891_ (.A(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__nor2_1 _12892_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_04030_),
    .Y(_05629_));
 sky130_fd_sc_hd__a31o_1 _12893_ (.A1(_04031_),
    .A2(_05329_),
    .A3(_05330_),
    .B1(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(_05454_),
    .A1(_05630_),
    .S(_05561_),
    .X(_05631_));
 sky130_fd_sc_hd__o211a_1 _12895_ (.A1(_05623_),
    .A2(_05626_),
    .B1(_05628_),
    .C1(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__o311a_1 _12896_ (.A1(_05609_),
    .A2(_05619_),
    .A3(_05622_),
    .B1(_05566_),
    .C1(_05562_),
    .X(_05633_));
 sky130_fd_sc_hd__xor2_2 _12897_ (.A(_05626_),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__o211a_1 _12898_ (.A1(_05609_),
    .A2(_05619_),
    .B1(_05562_),
    .C1(_05566_),
    .X(_05635_));
 sky130_fd_sc_hd__xor2_2 _12899_ (.A(_05622_),
    .B(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__a211o_1 _12900_ (.A1(_05628_),
    .A2(_05626_),
    .B1(_05633_),
    .C1(_05631_),
    .X(_05637_));
 sky130_fd_sc_hd__or4b_4 _12901_ (.A(_05632_),
    .B(_05634_),
    .C(_05636_),
    .D_N(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__and3_1 _12902_ (.A(_05562_),
    .B(_05566_),
    .C(_05601_),
    .X(_05639_));
 sky130_fd_sc_hd__xor2_2 _12903_ (.A(_05615_),
    .B(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__and3_1 _12904_ (.A(_05562_),
    .B(_05566_),
    .C(_05619_),
    .X(_05641_));
 sky130_fd_sc_hd__xor2_2 _12905_ (.A(_05609_),
    .B(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__a211o_1 _12906_ (.A1(_05610_),
    .A2(_05612_),
    .B1(_05615_),
    .C1(_05601_),
    .X(_05643_));
 sky130_fd_sc_hd__and3_1 _12907_ (.A(_05562_),
    .B(_05566_),
    .C(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__xor2_2 _12908_ (.A(_05618_),
    .B(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_2 _12909_ (.A(_05610_),
    .B(_05612_),
    .Y(_05646_));
 sky130_fd_sc_hd__o211a_1 _12910_ (.A1(_05615_),
    .A2(_05601_),
    .B1(_05566_),
    .C1(_05563_),
    .X(_05647_));
 sky130_fd_sc_hd__xnor2_4 _12911_ (.A(_05646_),
    .B(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__or4_2 _12912_ (.A(_05640_),
    .B(_05642_),
    .C(_05645_),
    .D(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__o41a_2 _12913_ (.A1(_05601_),
    .A2(_05606_),
    .A3(_05638_),
    .A4(_05649_),
    .B1(_05628_),
    .X(_05650_));
 sky130_fd_sc_hd__nor2_1 _12914_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_04031_),
    .Y(_05651_));
 sky130_fd_sc_hd__a211o_1 _12915_ (.A1(_04031_),
    .A2(_05372_),
    .B1(_05651_),
    .C1(_04001_),
    .X(_05652_));
 sky130_fd_sc_hd__a21o_1 _12916_ (.A1(\rbzero.wall_tracer.visualWallDist[7] ),
    .A2(_05571_),
    .B1(_05572_),
    .X(_05653_));
 sky130_fd_sc_hd__nand2_1 _12917_ (.A(_05563_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__a21oi_1 _12918_ (.A1(_05652_),
    .A2(_05654_),
    .B1(_05567_),
    .Y(_05655_));
 sky130_fd_sc_hd__nor2_1 _12919_ (.A(_05650_),
    .B(_05655_),
    .Y(_05656_));
 sky130_fd_sc_hd__o2111a_1 _12920_ (.A1(_05567_),
    .A2(_05575_),
    .B1(_05576_),
    .C1(_05656_),
    .D1(_05563_),
    .X(_05657_));
 sky130_fd_sc_hd__nor2_1 _12921_ (.A(_05567_),
    .B(_05576_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_1 _12922_ (.A(_04001_),
    .B(_05494_),
    .Y(_05659_));
 sky130_fd_sc_hd__and2_1 _12923_ (.A(_05659_),
    .B(_05569_),
    .X(_05660_));
 sky130_fd_sc_hd__nor2_1 _12924_ (.A(_05567_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__or3_1 _12925_ (.A(_05650_),
    .B(_05655_),
    .C(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__xnor2_1 _12926_ (.A(_05574_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__inv_2 _12927_ (.A(_05660_),
    .Y(_05664_));
 sky130_fd_sc_hd__or3_1 _12928_ (.A(_05650_),
    .B(_05655_),
    .C(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__o21ai_1 _12929_ (.A1(_05650_),
    .A2(_05655_),
    .B1(_05664_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_1 _12930_ (.A(_05652_),
    .B(_05659_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _12931_ (.A(_05628_),
    .B(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__o21bai_1 _12933_ (.A1(_05650_),
    .A2(_05669_),
    .B1_N(_05654_),
    .Y(_05670_));
 sky130_fd_sc_hd__a211o_1 _12934_ (.A1(_05563_),
    .A2(_05653_),
    .B1(_05669_),
    .C1(_05650_),
    .X(_05671_));
 sky130_fd_sc_hd__a22o_1 _12935_ (.A1(_05665_),
    .A2(_05666_),
    .B1(_05670_),
    .B2(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__or4_2 _12936_ (.A(_05657_),
    .B(_05658_),
    .C(_05663_),
    .D(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__xor2_1 _12937_ (.A(_05667_),
    .B(_05650_),
    .X(_05674_));
 sky130_fd_sc_hd__nand2_1 _12938_ (.A(_05659_),
    .B(_05603_),
    .Y(_05675_));
 sky130_fd_sc_hd__o41a_1 _12939_ (.A1(_05601_),
    .A2(_05604_),
    .A3(_05638_),
    .A4(_05649_),
    .B1(_05628_),
    .X(_05676_));
 sky130_fd_sc_hd__xor2_2 _12940_ (.A(_05675_),
    .B(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__clkinv_2 _12941_ (.A(_05605_),
    .Y(_05678_));
 sky130_fd_sc_hd__clkinv_2 _12942_ (.A(_05604_),
    .Y(_05679_));
 sky130_fd_sc_hd__o31a_1 _12943_ (.A1(_05601_),
    .A2(_05638_),
    .A3(_05649_),
    .B1(_05628_),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(_05678_),
    .A1(_05679_),
    .S(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__or2_1 _12945_ (.A(_05677_),
    .B(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__or2_2 _12946_ (.A(_05674_),
    .B(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__or2_2 _12947_ (.A(_05673_),
    .B(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__nand2_2 _12948_ (.A(_05577_),
    .B(_05579_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21a_1 _12949_ (.A1(_05582_),
    .A2(_05600_),
    .B1(_05628_),
    .X(_05686_));
 sky130_fd_sc_hd__xnor2_4 _12950_ (.A(_05685_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__inv_2 _12951_ (.A(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__or3_1 _12952_ (.A(_05638_),
    .B(_05649_),
    .C(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__or2b_2 _12953_ (.A(_05632_),
    .B_N(_05637_),
    .X(_05690_));
 sky130_fd_sc_hd__or2_1 _12954_ (.A(_05690_),
    .B(_05634_),
    .X(_05691_));
 sky130_fd_sc_hd__or2_1 _12955_ (.A(_05642_),
    .B(_05645_),
    .X(_05692_));
 sky130_fd_sc_hd__or3b_1 _12956_ (.A(_05692_),
    .B(_05636_),
    .C_N(_05648_),
    .X(_05693_));
 sky130_fd_sc_hd__or4_2 _12957_ (.A(_05691_),
    .B(_05673_),
    .C(_05683_),
    .D(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__buf_2 _12958_ (.A(_05674_),
    .X(_05695_));
 sky130_fd_sc_hd__or2_1 _12959_ (.A(_05638_),
    .B(_05682_),
    .X(_05696_));
 sky130_fd_sc_hd__xnor2_2 _12960_ (.A(_05615_),
    .B(_05639_),
    .Y(_05697_));
 sky130_fd_sc_hd__or3_1 _12961_ (.A(_05697_),
    .B(_05692_),
    .C(_05648_),
    .X(_05698_));
 sky130_fd_sc_hd__or4_2 _12962_ (.A(_05695_),
    .B(_05673_),
    .C(_05696_),
    .D(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__o211ai_4 _12963_ (.A1(_05684_),
    .A2(_05689_),
    .B1(_05694_),
    .C1(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__or3_2 _12964_ (.A(_05638_),
    .B(_05649_),
    .C(_05687_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_2 _12965_ (.A(_05673_),
    .X(_05702_));
 sky130_fd_sc_hd__nor3_4 _12966_ (.A(_05701_),
    .B(_05702_),
    .C(_05683_),
    .Y(_05703_));
 sky130_fd_sc_hd__o21a_1 _12967_ (.A1(_05591_),
    .A2(_05593_),
    .B1(_05628_),
    .X(_05704_));
 sky130_fd_sc_hd__xnor2_2 _12968_ (.A(_05589_),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__and3_1 _12969_ (.A(_05563_),
    .B(_05566_),
    .C(_05591_),
    .X(_05706_));
 sky130_fd_sc_hd__xnor2_1 _12970_ (.A(_05593_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_1 _12971_ (.A(_05591_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__and3_1 _12972_ (.A(_05563_),
    .B(_05566_),
    .C(_05600_),
    .X(_05709_));
 sky130_fd_sc_hd__xor2_4 _12973_ (.A(_05582_),
    .B(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__or2_2 _12974_ (.A(_05586_),
    .B(_05587_),
    .X(_05711_));
 sky130_fd_sc_hd__o41a_2 _12975_ (.A1(_05594_),
    .A2(_05596_),
    .A3(_05598_),
    .A4(_05584_),
    .B1(_05628_),
    .X(_05712_));
 sky130_fd_sc_hd__xor2_2 _12976_ (.A(_05711_),
    .B(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__nor2_2 _12977_ (.A(_05567_),
    .B(_05599_),
    .Y(_05714_));
 sky130_fd_sc_hd__xor2_2 _12978_ (.A(_05584_),
    .B(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__or3_1 _12979_ (.A(_05710_),
    .B(_05713_),
    .C(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__o21a_1 _12980_ (.A1(_05594_),
    .A2(_05596_),
    .B1(_05628_),
    .X(_05717_));
 sky130_fd_sc_hd__xor2_1 _12981_ (.A(_05598_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__or2_1 _12982_ (.A(_05716_),
    .B(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__and3_1 _12983_ (.A(_05563_),
    .B(_05566_),
    .C(_05594_),
    .X(_05720_));
 sky130_fd_sc_hd__xor2_4 _12984_ (.A(_05596_),
    .B(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__a211oi_1 _12985_ (.A1(_05705_),
    .A2(_05708_),
    .B1(_05719_),
    .C1(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__nand2_1 _12986_ (.A(_05670_),
    .B(_05671_),
    .Y(_05723_));
 sky130_fd_sc_hd__inv_2 _12987_ (.A(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _12988_ (.A(_05665_),
    .B(_05666_),
    .Y(_05725_));
 sky130_fd_sc_hd__or4b_1 _12989_ (.A(_05657_),
    .B(_05658_),
    .C(_05663_),
    .D_N(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__o21ba_1 _12990_ (.A1(_05724_),
    .A2(_05683_),
    .B1_N(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__xnor2_1 _12991_ (.A(_05609_),
    .B(_05641_),
    .Y(_05728_));
 sky130_fd_sc_hd__nand2_1 _12992_ (.A(_05728_),
    .B(_05645_),
    .Y(_05729_));
 sky130_fd_sc_hd__or4_1 _12993_ (.A(_05638_),
    .B(_05695_),
    .C(_05677_),
    .D(_05681_),
    .X(_05730_));
 sky130_fd_sc_hd__nor3_1 _12994_ (.A(_05702_),
    .B(_05729_),
    .C(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__a211o_1 _12995_ (.A1(_05703_),
    .A2(_05722_),
    .B1(_05727_),
    .C1(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__inv_2 _12996_ (.A(_05721_),
    .Y(_05733_));
 sky130_fd_sc_hd__xor2_2 _12997_ (.A(_05589_),
    .B(_05704_),
    .X(_05734_));
 sky130_fd_sc_hd__or3_1 _12998_ (.A(_05721_),
    .B(_05734_),
    .C(_05707_),
    .X(_05735_));
 sky130_fd_sc_hd__or2_2 _12999_ (.A(_05687_),
    .B(_05719_),
    .X(_05736_));
 sky130_fd_sc_hd__or4_4 _13000_ (.A(_05649_),
    .B(_05695_),
    .C(_05673_),
    .D(_05696_),
    .X(_05737_));
 sky130_fd_sc_hd__a211o_1 _13001_ (.A1(_05733_),
    .A2(_05735_),
    .B1(_05736_),
    .C1(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__or3b_1 _13002_ (.A(_05700_),
    .B(_05732_),
    .C_N(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__clkbuf_2 _13003_ (.A(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__buf_2 _13004_ (.A(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__clkbuf_4 _13005_ (.A(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__nor3b_2 _13006_ (.A(_05700_),
    .B(_05732_),
    .C_N(_05738_),
    .Y(_05743_));
 sky130_fd_sc_hd__xnor2_2 _13007_ (.A(_05622_),
    .B(_05635_),
    .Y(_05744_));
 sky130_fd_sc_hd__a21oi_1 _13008_ (.A1(_05642_),
    .A2(_05744_),
    .B1(_05634_),
    .Y(_05745_));
 sky130_fd_sc_hd__or4_1 _13009_ (.A(_05690_),
    .B(_05702_),
    .C(_05683_),
    .D(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__inv_2 _13010_ (.A(_05690_),
    .Y(_05747_));
 sky130_fd_sc_hd__or3_1 _13011_ (.A(_05691_),
    .B(_05744_),
    .C(_05682_),
    .X(_05748_));
 sky130_fd_sc_hd__or3_1 _13012_ (.A(_05695_),
    .B(_05702_),
    .C(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__or3_1 _13013_ (.A(_05601_),
    .B(_05638_),
    .C(_05649_),
    .X(_05750_));
 sky130_fd_sc_hd__or3_1 _13014_ (.A(_05750_),
    .B(_05702_),
    .C(_05683_),
    .X(_05751_));
 sky130_fd_sc_hd__buf_4 _13015_ (.A(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__o211a_1 _13016_ (.A1(_05747_),
    .A2(_05684_),
    .B1(_05749_),
    .C1(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__and4bb_2 _13017_ (.A_N(_05700_),
    .B_N(_05731_),
    .C(_05746_),
    .D(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__or2_1 _13018_ (.A(_05743_),
    .B(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__or2_1 _13019_ (.A(_05736_),
    .B(_05735_),
    .X(_05756_));
 sky130_fd_sc_hd__xnor2_2 _13020_ (.A(_05584_),
    .B(_05714_),
    .Y(_05757_));
 sky130_fd_sc_hd__or4_1 _13021_ (.A(_05710_),
    .B(_05713_),
    .C(_05757_),
    .D(_05687_),
    .X(_05758_));
 sky130_fd_sc_hd__a21oi_1 _13022_ (.A1(_05756_),
    .A2(_05758_),
    .B1(_05737_),
    .Y(_05759_));
 sky130_fd_sc_hd__or2_1 _13023_ (.A(_05695_),
    .B(_05702_),
    .X(_05760_));
 sky130_fd_sc_hd__inv_2 _13024_ (.A(_05677_),
    .Y(_05761_));
 sky130_fd_sc_hd__mux2_1 _13025_ (.A0(_05605_),
    .A1(_05604_),
    .S(_05680_),
    .X(_05762_));
 sky130_fd_sc_hd__and3_1 _13026_ (.A(_05761_),
    .B(_05762_),
    .C(_05748_),
    .X(_05763_));
 sky130_fd_sc_hd__xor2_1 _13027_ (.A(_05574_),
    .B(_05662_),
    .X(_05764_));
 sky130_fd_sc_hd__o21a_1 _13028_ (.A1(_05567_),
    .A2(_05575_),
    .B1(_05656_),
    .X(_05765_));
 sky130_fd_sc_hd__o21ba_1 _13029_ (.A1(_05765_),
    .A2(_05576_),
    .B1_N(_05657_),
    .X(_05766_));
 sky130_fd_sc_hd__a21bo_1 _13030_ (.A1(_05725_),
    .A2(_05764_),
    .B1_N(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__nand2_1 _13031_ (.A(_05642_),
    .B(_05744_),
    .Y(_05768_));
 sky130_fd_sc_hd__or4_1 _13032_ (.A(_05691_),
    .B(_05673_),
    .C(_05683_),
    .D(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__or4_1 _13033_ (.A(_05719_),
    .B(_05721_),
    .C(_05734_),
    .D(_05708_),
    .X(_05770_));
 sky130_fd_sc_hd__or4_1 _13034_ (.A(_05701_),
    .B(_05702_),
    .C(_05683_),
    .D(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__o2111ai_2 _13035_ (.A1(_05760_),
    .A2(_05763_),
    .B1(_05767_),
    .C1(_05769_),
    .D1(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__xnor2_2 _13036_ (.A(_05598_),
    .B(_05717_),
    .Y(_05773_));
 sky130_fd_sc_hd__nor2_1 _13037_ (.A(_05716_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__a2bb2o_2 _13038_ (.A1_N(_05684_),
    .A2_N(_05689_),
    .B1(_05703_),
    .B2(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__or4b_1 _13039_ (.A(_05759_),
    .B(_05772_),
    .C(_05775_),
    .D_N(_05699_),
    .X(_05776_));
 sky130_fd_sc_hd__clkbuf_2 _13040_ (.A(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__clkbuf_4 _13041_ (.A(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__buf_2 _13042_ (.A(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__or4_1 _13043_ (.A(_05695_),
    .B(_05702_),
    .C(_05677_),
    .D(_05762_),
    .X(_05780_));
 sky130_fd_sc_hd__clkinv_2 _13044_ (.A(_05695_),
    .Y(_05781_));
 sky130_fd_sc_hd__or2_1 _13045_ (.A(_05781_),
    .B(_05702_),
    .X(_05782_));
 sky130_fd_sc_hd__xnor2_2 _13046_ (.A(_05711_),
    .B(_05712_),
    .Y(_05783_));
 sky130_fd_sc_hd__o32a_1 _13047_ (.A1(_05719_),
    .A2(_05721_),
    .A3(_05705_),
    .B1(_05783_),
    .B2(_05710_),
    .X(_05784_));
 sky130_fd_sc_hd__or3_1 _13048_ (.A(_05701_),
    .B(_05682_),
    .C(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__or4_1 _13049_ (.A(_05725_),
    .B(_05657_),
    .C(_05658_),
    .D(_05663_),
    .X(_05786_));
 sky130_fd_sc_hd__o311a_1 _13050_ (.A1(_05695_),
    .A2(_05702_),
    .A3(_05785_),
    .B1(_05786_),
    .C1(_05766_),
    .X(_05787_));
 sky130_fd_sc_hd__nand4_2 _13051_ (.A(_05780_),
    .B(_05746_),
    .C(_05782_),
    .D(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__nand2_1 _13052_ (.A(_05694_),
    .B(_05771_),
    .Y(_05789_));
 sky130_fd_sc_hd__or3_1 _13053_ (.A(_05775_),
    .B(_05788_),
    .C(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__clkbuf_4 _13054_ (.A(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_4 _13055_ (.A(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__clkbuf_4 _13056_ (.A(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__inv_2 _13057_ (.A(_05700_),
    .Y(_05794_));
 sky130_fd_sc_hd__nor4b_2 _13058_ (.A(_05759_),
    .B(_05772_),
    .C(_05775_),
    .D_N(_05699_),
    .Y(_05795_));
 sky130_fd_sc_hd__nor3_4 _13059_ (.A(_05775_),
    .B(_05788_),
    .C(_05789_),
    .Y(_05796_));
 sky130_fd_sc_hd__a21o_1 _13060_ (.A1(_05795_),
    .A2(_05796_),
    .B1(_05743_),
    .X(_05797_));
 sky130_fd_sc_hd__nand2_2 _13061_ (.A(_05754_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _13062_ (.A(_05794_),
    .B(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__buf_4 _13063_ (.A(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__clkbuf_4 _13064_ (.A(_05796_),
    .X(_05801_));
 sky130_fd_sc_hd__mux4_1 _13065_ (.A0(_05710_),
    .A1(_05715_),
    .A2(_05718_),
    .A3(_05713_),
    .S0(_05777_),
    .S1(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__xor2_2 _13066_ (.A(_05593_),
    .B(_05706_),
    .X(_05803_));
 sky130_fd_sc_hd__mux2_1 _13067_ (.A0(_05591_),
    .A1(_05803_),
    .S(_05791_),
    .X(_05804_));
 sky130_fd_sc_hd__mux2_1 _13068_ (.A0(_05721_),
    .A1(_05734_),
    .S(_05796_),
    .X(_05805_));
 sky130_fd_sc_hd__xnor2_1 _13069_ (.A(_05777_),
    .B(_05796_),
    .Y(_05806_));
 sky130_fd_sc_hd__clkbuf_4 _13070_ (.A(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__mux2_1 _13071_ (.A0(_05804_),
    .A1(_05805_),
    .S(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__or3_1 _13072_ (.A(_05740_),
    .B(_05777_),
    .C(_05790_),
    .X(_05809_));
 sky130_fd_sc_hd__and2_1 _13073_ (.A(_05797_),
    .B(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__buf_2 _13074_ (.A(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _13075_ (.A0(_05802_),
    .A1(_05808_),
    .S(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__a21oi_1 _13076_ (.A1(_05754_),
    .A2(_05797_),
    .B1(_05700_),
    .Y(_05813_));
 sky130_fd_sc_hd__clkbuf_4 _13077_ (.A(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__mux4_1 _13078_ (.A0(_05640_),
    .A1(_05645_),
    .A2(_05648_),
    .A3(_05687_),
    .S0(_05795_),
    .S1(_05801_),
    .X(_05815_));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(_05642_),
    .A1(_05636_),
    .S(_05791_),
    .X(_05816_));
 sky130_fd_sc_hd__or4_1 _13080_ (.A(_05634_),
    .B(_05775_),
    .C(_05788_),
    .D(_05789_),
    .X(_05817_));
 sky130_fd_sc_hd__o21a_1 _13081_ (.A1(_05690_),
    .A2(_05796_),
    .B1(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__mux2_1 _13082_ (.A0(_05816_),
    .A1(_05818_),
    .S(_05806_),
    .X(_05819_));
 sky130_fd_sc_hd__nand2_2 _13083_ (.A(_05797_),
    .B(_05809_),
    .Y(_05820_));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(_05815_),
    .A1(_05819_),
    .S(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__or2_1 _13085_ (.A(_05814_),
    .B(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__o21ai_4 _13086_ (.A1(_05800_),
    .A2(_05812_),
    .B1(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__clkbuf_4 _13087_ (.A(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__buf_4 _13088_ (.A(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_4 _13089_ (.A(_05795_),
    .X(_05826_));
 sky130_fd_sc_hd__mux2_1 _13090_ (.A0(_05591_),
    .A1(_05803_),
    .S(_05796_),
    .X(_05827_));
 sky130_fd_sc_hd__and2_1 _13091_ (.A(_05826_),
    .B(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__mux2_1 _13092_ (.A0(_05757_),
    .A1(_05773_),
    .S(_05792_),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _13093_ (.A0(_05733_),
    .A1(_05705_),
    .S(_05792_),
    .X(_05830_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(_05829_),
    .A1(_05830_),
    .S(_05778_),
    .X(_05831_));
 sky130_fd_sc_hd__nand2_1 _13095_ (.A(_05740_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__or2_1 _13096_ (.A(_05700_),
    .B(_05703_),
    .X(_05833_));
 sky130_fd_sc_hd__clkbuf_4 _13097_ (.A(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__o211a_1 _13098_ (.A1(_05740_),
    .A2(_05828_),
    .B1(_05832_),
    .C1(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__mux2_1 _13099_ (.A0(_05640_),
    .A1(_05648_),
    .S(_05791_),
    .X(_05836_));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(_05642_),
    .A1(_05645_),
    .S(_05796_),
    .X(_05837_));
 sky130_fd_sc_hd__mux2_1 _13101_ (.A0(_05836_),
    .A1(_05837_),
    .S(_05807_),
    .X(_05838_));
 sky130_fd_sc_hd__mux4_1 _13102_ (.A0(_05710_),
    .A1(_05713_),
    .A2(_05715_),
    .A3(_05687_),
    .S0(_05791_),
    .S1(_05826_),
    .X(_05839_));
 sky130_fd_sc_hd__mux2_1 _13103_ (.A0(_05838_),
    .A1(_05839_),
    .S(_05811_),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(_05634_),
    .A1(_05636_),
    .S(_05796_),
    .X(_05841_));
 sky130_fd_sc_hd__mux2_1 _13105_ (.A0(_05690_),
    .A1(_05681_),
    .S(_05791_),
    .X(_05842_));
 sky130_fd_sc_hd__mux2_1 _13106_ (.A0(_05841_),
    .A1(_05842_),
    .S(_05807_),
    .X(_05843_));
 sky130_fd_sc_hd__clkbuf_4 _13107_ (.A(_05811_),
    .X(_05844_));
 sky130_fd_sc_hd__a22o_1 _13108_ (.A1(_05814_),
    .A2(_05840_),
    .B1(_05843_),
    .B2(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__nor2_4 _13109_ (.A(_05835_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(_05798_),
    .Y(_05847_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(_05838_),
    .A1(_05843_),
    .S(_05820_),
    .X(_05848_));
 sky130_fd_sc_hd__mux4_1 _13112_ (.A0(_05718_),
    .A1(_05734_),
    .A2(_05803_),
    .A3(_05721_),
    .S0(_05777_),
    .S1(_05801_),
    .X(_05849_));
 sky130_fd_sc_hd__a21o_1 _13113_ (.A1(_05797_),
    .A2(_05809_),
    .B1(_05839_),
    .X(_05850_));
 sky130_fd_sc_hd__o211a_1 _13114_ (.A1(_05820_),
    .A2(_05849_),
    .B1(_05850_),
    .C1(_05798_),
    .X(_05851_));
 sky130_fd_sc_hd__a211o_2 _13115_ (.A1(_05847_),
    .A2(_05848_),
    .B1(_05851_),
    .C1(_05700_),
    .X(_05852_));
 sky130_fd_sc_hd__or2_2 _13116_ (.A(_05794_),
    .B(_05828_),
    .X(_05853_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(_05812_),
    .A1(_05821_),
    .S(_05799_),
    .X(_05854_));
 sky130_fd_sc_hd__clkbuf_4 _13118_ (.A(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__a21o_1 _13119_ (.A1(_05852_),
    .A2(_05853_),
    .B1(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__o21ai_1 _13120_ (.A1(_05690_),
    .A2(_05801_),
    .B1(_05817_),
    .Y(_05857_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(_05761_),
    .A1(_05762_),
    .S(_05796_),
    .X(_05858_));
 sky130_fd_sc_hd__mux2_1 _13122_ (.A0(_05857_),
    .A1(_05858_),
    .S(_05807_),
    .X(_05859_));
 sky130_fd_sc_hd__or4_1 _13123_ (.A(_05648_),
    .B(_05775_),
    .C(_05788_),
    .D(_05789_),
    .X(_05860_));
 sky130_fd_sc_hd__o21ai_1 _13124_ (.A1(_05645_),
    .A2(_05796_),
    .B1(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(_05728_),
    .A1(_05744_),
    .S(_05791_),
    .X(_05862_));
 sky130_fd_sc_hd__mux2_1 _13126_ (.A0(_05861_),
    .A1(_05862_),
    .S(_05807_),
    .X(_05863_));
 sky130_fd_sc_hd__mux2_1 _13127_ (.A0(_05859_),
    .A1(_05863_),
    .S(_05811_),
    .X(_05864_));
 sky130_fd_sc_hd__nor2_1 _13128_ (.A(_05798_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__mux4_1 _13129_ (.A0(_05715_),
    .A1(_05721_),
    .A2(_05734_),
    .A3(_05718_),
    .S0(_05777_),
    .S1(_05801_),
    .X(_05866_));
 sky130_fd_sc_hd__inv_2 _13130_ (.A(_05710_),
    .Y(_05867_));
 sky130_fd_sc_hd__mux4_1 _13131_ (.A0(_05867_),
    .A1(_05697_),
    .A2(_05688_),
    .A3(_05783_),
    .S0(_05826_),
    .S1(_05801_),
    .X(_05868_));
 sky130_fd_sc_hd__nand2_1 _13132_ (.A(_05820_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__o211a_1 _13133_ (.A1(_05820_),
    .A2(_05866_),
    .B1(_05869_),
    .C1(_05813_),
    .X(_05870_));
 sky130_fd_sc_hd__nor2_2 _13134_ (.A(_05700_),
    .B(_05703_),
    .Y(_05871_));
 sky130_fd_sc_hd__mux2_1 _13135_ (.A0(_05705_),
    .A1(_05707_),
    .S(_05791_),
    .X(_05872_));
 sky130_fd_sc_hd__or3b_1 _13136_ (.A(_05791_),
    .B(_05795_),
    .C_N(_05591_),
    .X(_05873_));
 sky130_fd_sc_hd__o21a_1 _13137_ (.A1(_05778_),
    .A2(_05872_),
    .B1(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__or3_1 _13138_ (.A(_05703_),
    .B(_05871_),
    .C(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__or3b_1 _13139_ (.A(_05865_),
    .B(_05870_),
    .C_N(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__buf_2 _13140_ (.A(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__clkinv_2 _13141_ (.A(_05827_),
    .Y(_05878_));
 sky130_fd_sc_hd__mux2_2 _13142_ (.A0(_05830_),
    .A1(_05878_),
    .S(_05778_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_1 _13143_ (.A0(_05837_),
    .A1(_05841_),
    .S(_05807_),
    .X(_05880_));
 sky130_fd_sc_hd__a21oi_2 _13144_ (.A1(_05844_),
    .A2(_05880_),
    .B1(_05798_),
    .Y(_05881_));
 sky130_fd_sc_hd__mux4_1 _13145_ (.A0(_05710_),
    .A1(_05640_),
    .A2(_05648_),
    .A3(_05687_),
    .S0(_05778_),
    .S1(_05792_),
    .X(_05882_));
 sky130_fd_sc_hd__nor2_1 _13146_ (.A(_05844_),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__clkbuf_4 _13147_ (.A(_05820_),
    .X(_05884_));
 sky130_fd_sc_hd__mux4_1 _13148_ (.A0(_05713_),
    .A1(_05718_),
    .A2(_05721_),
    .A3(_05715_),
    .S0(_05778_),
    .S1(_05801_),
    .X(_05885_));
 sky130_fd_sc_hd__nor2_1 _13149_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__o21a_1 _13150_ (.A1(_05883_),
    .A2(_05886_),
    .B1(_05798_),
    .X(_05887_));
 sky130_fd_sc_hd__a211oi_4 _13151_ (.A1(_05700_),
    .A2(_05879_),
    .B1(_05881_),
    .C1(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__a21o_2 _13152_ (.A1(_05856_),
    .A2(_05877_),
    .B1(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(_05773_),
    .A1(_05733_),
    .S(_05792_),
    .X(_05890_));
 sky130_fd_sc_hd__mux2_1 _13154_ (.A0(_05872_),
    .A1(_05890_),
    .S(_05826_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_4 _13155_ (.A(_05743_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_4 _13156_ (.A(_05801_),
    .X(_05893_));
 sky130_fd_sc_hd__and3_1 _13157_ (.A(_05743_),
    .B(_05826_),
    .C(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__a2bb2o_1 _13158_ (.A1_N(_05891_),
    .A2_N(_05892_),
    .B1(_05591_),
    .B2(_05894_),
    .X(_05895_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(_05802_),
    .A1(_05815_),
    .S(_05884_),
    .X(_05896_));
 sky130_fd_sc_hd__a21o_1 _13160_ (.A1(_05811_),
    .A2(_05819_),
    .B1(_05814_),
    .X(_05897_));
 sky130_fd_sc_hd__o21a_1 _13161_ (.A1(_05800_),
    .A2(_05896_),
    .B1(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__a21oi_4 _13162_ (.A1(_05834_),
    .A2(_05895_),
    .B1(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__nor2_1 _13163_ (.A(_05846_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__and2_2 _13164_ (.A(_05743_),
    .B(_05754_),
    .X(_05901_));
 sky130_fd_sc_hd__inv_2 _13165_ (.A(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(_05783_),
    .A1(_05757_),
    .S(_05791_),
    .X(_05903_));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(_05890_),
    .A1(_05903_),
    .S(_05826_),
    .X(_05904_));
 sky130_fd_sc_hd__o22a_1 _13168_ (.A1(_05902_),
    .A2(_05874_),
    .B1(_05904_),
    .B2(_05755_),
    .X(_05905_));
 sky130_fd_sc_hd__mux2_1 _13169_ (.A0(_05863_),
    .A1(_05868_),
    .S(_05811_),
    .X(_05906_));
 sky130_fd_sc_hd__or2_1 _13170_ (.A(_05800_),
    .B(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__or2_1 _13171_ (.A(_05884_),
    .B(_05859_),
    .X(_05908_));
 sky130_fd_sc_hd__o211a_2 _13172_ (.A1(_05871_),
    .A2(_05905_),
    .B1(_05907_),
    .C1(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__inv_2 _13173_ (.A(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(_05867_),
    .A1(_05783_),
    .S(_05792_),
    .X(_05911_));
 sky130_fd_sc_hd__a21o_1 _13175_ (.A1(_05826_),
    .A2(_05911_),
    .B1(_05755_),
    .X(_05912_));
 sky130_fd_sc_hd__a21o_1 _13176_ (.A1(_05778_),
    .A2(_05829_),
    .B1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__or2_1 _13177_ (.A(_05902_),
    .B(_05879_),
    .X(_05914_));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(_05880_),
    .A1(_05882_),
    .S(_05811_),
    .X(_05915_));
 sky130_fd_sc_hd__mux2_1 _13179_ (.A0(_05695_),
    .A1(_05677_),
    .S(_05801_),
    .X(_05916_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(_05842_),
    .A1(_05916_),
    .S(_05807_),
    .X(_05917_));
 sky130_fd_sc_hd__a21o_1 _13181_ (.A1(_05844_),
    .A2(_05917_),
    .B1(_05834_),
    .X(_05918_));
 sky130_fd_sc_hd__a21oi_1 _13182_ (.A1(_05814_),
    .A2(_05915_),
    .B1(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__a31o_2 _13183_ (.A1(_05834_),
    .A2(_05913_),
    .A3(_05914_),
    .B1(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__clkinv_2 _13184_ (.A(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__a31o_1 _13185_ (.A1(_05889_),
    .A2(_05900_),
    .A3(_05910_),
    .B1(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__buf_4 _13186_ (.A(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__mux2_1 _13187_ (.A0(_05695_),
    .A1(_05724_),
    .S(_05793_),
    .X(_05924_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_05807_),
    .B(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__o21ai_1 _13189_ (.A1(_05807_),
    .A2(_05858_),
    .B1(_05871_),
    .Y(_05926_));
 sky130_fd_sc_hd__a21oi_1 _13190_ (.A1(_05814_),
    .A2(_05821_),
    .B1(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__nor2_2 _13191_ (.A(_05743_),
    .B(_05754_),
    .Y(_05928_));
 sky130_fd_sc_hd__nor2_2 _13192_ (.A(_05703_),
    .B(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__a21oi_1 _13193_ (.A1(_05901_),
    .A2(_05891_),
    .B1(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__buf_2 _13194_ (.A(_05826_),
    .X(_05931_));
 sky130_fd_sc_hd__or2_1 _13195_ (.A(_05928_),
    .B(_05901_),
    .X(_05932_));
 sky130_fd_sc_hd__a41o_1 _13196_ (.A1(_05591_),
    .A2(_05740_),
    .A3(_05931_),
    .A4(_05893_),
    .B1(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__mux2_1 _13197_ (.A0(_05867_),
    .A1(_05688_),
    .S(_05801_),
    .X(_05934_));
 sky130_fd_sc_hd__o21a_1 _13198_ (.A1(_05778_),
    .A2(_05934_),
    .B1(_05928_),
    .X(_05935_));
 sky130_fd_sc_hd__o21ai_1 _13199_ (.A1(_05931_),
    .A2(_05903_),
    .B1(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__a31o_1 _13200_ (.A1(_05930_),
    .A2(_05933_),
    .A3(_05936_),
    .B1(_05871_),
    .X(_05937_));
 sky130_fd_sc_hd__a21bo_1 _13201_ (.A1(_05925_),
    .A2(_05927_),
    .B1_N(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__buf_4 _13202_ (.A(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__xnor2_4 _13203_ (.A(_05923_),
    .B(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_1 _13204_ (.A(_05889_),
    .B(_05900_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_1 _13205_ (.A1(_05941_),
    .A2(_05910_),
    .B1(_05923_),
    .Y(_05942_));
 sky130_fd_sc_hd__or3_1 _13206_ (.A(_05846_),
    .B(_05940_),
    .C(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__a211o_1 _13207_ (.A1(_05700_),
    .A2(_05879_),
    .B1(_05881_),
    .C1(_05887_),
    .X(_05944_));
 sky130_fd_sc_hd__a21o_2 _13208_ (.A1(_05856_),
    .A2(_05877_),
    .B1(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__a21oi_2 _13209_ (.A1(_05852_),
    .A2(_05853_),
    .B1(_05855_),
    .Y(_05946_));
 sky130_fd_sc_hd__nor3b_1 _13210_ (.A(_05865_),
    .B(_05870_),
    .C_N(_05875_),
    .Y(_05947_));
 sky130_fd_sc_hd__or3_1 _13211_ (.A(_05946_),
    .B(_05947_),
    .C(_05888_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_2 _13212_ (.A(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__inv_2 _13213_ (.A(_05848_),
    .Y(_05950_));
 sky130_fd_sc_hd__xnor2_1 _13214_ (.A(_05826_),
    .B(_05893_),
    .Y(_05951_));
 sky130_fd_sc_hd__clkbuf_4 _13215_ (.A(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__mux2_1 _13216_ (.A0(_05725_),
    .A1(_05723_),
    .S(_05893_),
    .X(_05953_));
 sky130_fd_sc_hd__nor2_1 _13217_ (.A(_05952_),
    .B(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__a21oi_1 _13218_ (.A1(_05952_),
    .A2(_05916_),
    .B1(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__a21oi_1 _13219_ (.A1(_05740_),
    .A2(_05828_),
    .B1(_05932_),
    .Y(_05956_));
 sky130_fd_sc_hd__nor2_1 _13220_ (.A(_05640_),
    .B(_05792_),
    .Y(_05957_));
 sky130_fd_sc_hd__a211o_1 _13221_ (.A1(_05688_),
    .A2(_05792_),
    .B1(_05957_),
    .C1(_05778_),
    .X(_05958_));
 sky130_fd_sc_hd__o211a_1 _13222_ (.A1(_05931_),
    .A2(_05911_),
    .B1(_05958_),
    .C1(_05928_),
    .X(_05959_));
 sky130_fd_sc_hd__a2111o_1 _13223_ (.A1(_05901_),
    .A2(_05831_),
    .B1(_05956_),
    .C1(_05959_),
    .D1(_05871_),
    .X(_05960_));
 sky130_fd_sc_hd__o211a_2 _13224_ (.A1(_05800_),
    .A2(_05950_),
    .B1(_05955_),
    .C1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__a21oi_2 _13225_ (.A1(_05945_),
    .A2(_05949_),
    .B1(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__nor2_1 _13226_ (.A(_05928_),
    .B(_05901_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21a_1 _13227_ (.A1(_05743_),
    .A2(_05874_),
    .B1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__a21o_1 _13228_ (.A1(_05697_),
    .A2(_05792_),
    .B1(_05778_),
    .X(_05965_));
 sky130_fd_sc_hd__nor2_1 _13229_ (.A(_05648_),
    .B(_05792_),
    .Y(_05966_));
 sky130_fd_sc_hd__o221a_1 _13230_ (.A1(_05826_),
    .A2(_05934_),
    .B1(_05965_),
    .B2(_05966_),
    .C1(_05928_),
    .X(_05967_));
 sky130_fd_sc_hd__or2_1 _13231_ (.A(_05929_),
    .B(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__a211o_1 _13232_ (.A1(_05901_),
    .A2(_05904_),
    .B1(_05964_),
    .C1(_05968_),
    .X(_05969_));
 sky130_fd_sc_hd__nand2_1 _13233_ (.A(_05951_),
    .B(_05924_),
    .Y(_05970_));
 sky130_fd_sc_hd__mux2_1 _13234_ (.A0(_05725_),
    .A1(_05764_),
    .S(_05793_),
    .X(_05971_));
 sky130_fd_sc_hd__o211a_1 _13235_ (.A1(_05800_),
    .A2(_05864_),
    .B1(_05970_),
    .C1(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__mux2_2 _13236_ (.A0(_05969_),
    .A1(_05972_),
    .S(_05871_),
    .X(_05973_));
 sky130_fd_sc_hd__buf_2 _13237_ (.A(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__xnor2_4 _13238_ (.A(_05889_),
    .B(_05899_),
    .Y(_05975_));
 sky130_fd_sc_hd__nor2_2 _13239_ (.A(_05974_),
    .B(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__nand2_1 _13240_ (.A(_05962_),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__buf_2 _13241_ (.A(_05939_),
    .X(_05978_));
 sky130_fd_sc_hd__a21oi_1 _13242_ (.A1(_05856_),
    .A2(_05877_),
    .B1(_05888_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21ai_2 _13243_ (.A1(_05979_),
    .A2(_05899_),
    .B1(_05846_),
    .Y(_05980_));
 sky130_fd_sc_hd__and2_1 _13244_ (.A(_05941_),
    .B(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__clkbuf_4 _13245_ (.A(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__buf_2 _13246_ (.A(_05961_),
    .X(_05983_));
 sky130_fd_sc_hd__and2_2 _13247_ (.A(_05945_),
    .B(_05949_),
    .X(_05984_));
 sky130_fd_sc_hd__o22a_1 _13248_ (.A1(_05983_),
    .A2(_05975_),
    .B1(_05984_),
    .B2(_05974_),
    .X(_05985_));
 sky130_fd_sc_hd__a21o_1 _13249_ (.A1(_05962_),
    .A2(_05976_),
    .B1(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__or3_1 _13250_ (.A(_05978_),
    .B(_05982_),
    .C(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_4 _13251_ (.A(_05941_),
    .X(_05988_));
 sky130_fd_sc_hd__clkinv_2 _13252_ (.A(_05939_),
    .Y(_05989_));
 sky130_fd_sc_hd__clkbuf_4 _13253_ (.A(_05909_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_4 _13254_ (.A(_05920_),
    .X(_05991_));
 sky130_fd_sc_hd__nand2_1 _13255_ (.A(_05990_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__and3_1 _13256_ (.A(_05988_),
    .B(_05989_),
    .C(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__or3b_1 _13257_ (.A(_05979_),
    .B(_05909_),
    .C_N(_05900_),
    .X(_05994_));
 sky130_fd_sc_hd__buf_2 _13258_ (.A(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__a22o_1 _13259_ (.A1(_05988_),
    .A2(_05989_),
    .B1(_05992_),
    .B2(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__or2b_1 _13260_ (.A(_05993_),
    .B_N(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__a21oi_1 _13261_ (.A1(_05977_),
    .A2(_05987_),
    .B1(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__and3_1 _13262_ (.A(_05977_),
    .B(_05987_),
    .C(_05997_),
    .X(_05999_));
 sky130_fd_sc_hd__nor2_1 _13263_ (.A(_05998_),
    .B(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__xnor2_1 _13264_ (.A(_05943_),
    .B(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__nand2_4 _13265_ (.A(_05945_),
    .B(_05949_),
    .Y(_06002_));
 sky130_fd_sc_hd__xnor2_1 _13266_ (.A(_06002_),
    .B(_05976_),
    .Y(_06003_));
 sky130_fd_sc_hd__or3_1 _13267_ (.A(_05983_),
    .B(_05981_),
    .C(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__o21ai_1 _13268_ (.A1(_05983_),
    .A2(_05982_),
    .B1(_06003_),
    .Y(_06005_));
 sky130_fd_sc_hd__nand2_1 _13269_ (.A(_06004_),
    .B(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__and3_1 _13270_ (.A(_05852_),
    .B(_05853_),
    .C(_05855_),
    .X(_06007_));
 sky130_fd_sc_hd__or2_1 _13271_ (.A(_05946_),
    .B(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_4 _13272_ (.A(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__nor2_1 _13273_ (.A(_05973_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__xnor2_1 _13274_ (.A(_05946_),
    .B(_05877_),
    .Y(_06011_));
 sky130_fd_sc_hd__inv_2 _13275_ (.A(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__nor2_1 _13276_ (.A(_05978_),
    .B(_05981_),
    .Y(_06013_));
 sky130_fd_sc_hd__xnor2_2 _13277_ (.A(_05986_),
    .B(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__nor2_2 _13278_ (.A(_05750_),
    .B(_05684_),
    .Y(_06015_));
 sky130_fd_sc_hd__clkbuf_4 _13279_ (.A(_06011_),
    .X(_06016_));
 sky130_fd_sc_hd__or2_1 _13280_ (.A(_06015_),
    .B(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__nor2_1 _13281_ (.A(_06010_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__a22o_1 _13282_ (.A1(_06010_),
    .A2(_06012_),
    .B1(_06014_),
    .B2(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__xnor2_1 _13283_ (.A(_06006_),
    .B(_06019_),
    .Y(_06020_));
 sky130_fd_sc_hd__xnor2_1 _13284_ (.A(_06001_),
    .B(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__xor2_2 _13285_ (.A(_06014_),
    .B(_06018_),
    .X(_06022_));
 sky130_fd_sc_hd__o21a_1 _13286_ (.A1(_05973_),
    .A2(_06011_),
    .B1(_06009_),
    .X(_06023_));
 sky130_fd_sc_hd__a21o_1 _13287_ (.A1(_06010_),
    .A2(_06012_),
    .B1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__nor2_1 _13288_ (.A(_05983_),
    .B(_06016_),
    .Y(_06025_));
 sky130_fd_sc_hd__or3_1 _13289_ (.A(_05946_),
    .B(_05973_),
    .C(_06007_),
    .X(_06026_));
 sky130_fd_sc_hd__xnor2_1 _13290_ (.A(_05855_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__a22o_1 _13291_ (.A1(_05855_),
    .A2(_06010_),
    .B1(_06025_),
    .B2(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__inv_2 _13292_ (.A(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__xor2_1 _13293_ (.A(_06024_),
    .B(_06028_),
    .X(_06030_));
 sky130_fd_sc_hd__clkbuf_4 _13294_ (.A(_05975_),
    .X(_06031_));
 sky130_fd_sc_hd__o21bai_1 _13295_ (.A1(_05978_),
    .A2(_06031_),
    .B1_N(_05962_),
    .Y(_06032_));
 sky130_fd_sc_hd__or3b_1 _13296_ (.A(_05939_),
    .B(_05975_),
    .C_N(_05962_),
    .X(_06033_));
 sky130_fd_sc_hd__a21oi_1 _13297_ (.A1(_05988_),
    .A2(_05980_),
    .B1(_05991_),
    .Y(_06034_));
 sky130_fd_sc_hd__a21o_1 _13298_ (.A1(_06032_),
    .A2(_06033_),
    .B1(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__nand3_1 _13299_ (.A(_06032_),
    .B(_06033_),
    .C(_06034_),
    .Y(_06036_));
 sky130_fd_sc_hd__nand3b_1 _13300_ (.A_N(_06030_),
    .B(_06035_),
    .C(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__o21ai_2 _13301_ (.A1(_06024_),
    .A2(_06029_),
    .B1(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__xnor2_1 _13302_ (.A(_06022_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_1 _13303_ (.A(_06033_),
    .B(_06036_),
    .Y(_06040_));
 sky130_fd_sc_hd__buf_2 _13304_ (.A(_05846_),
    .X(_06041_));
 sky130_fd_sc_hd__o21ai_1 _13305_ (.A1(_06041_),
    .A2(_05940_),
    .B1(_05942_),
    .Y(_06042_));
 sky130_fd_sc_hd__and2_1 _13306_ (.A(_05943_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__xnor2_1 _13307_ (.A(_06040_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__clkbuf_4 _13308_ (.A(_05899_),
    .X(_06045_));
 sky130_fd_sc_hd__or4_1 _13309_ (.A(_06041_),
    .B(_06045_),
    .C(_05991_),
    .D(_05978_),
    .X(_06046_));
 sky130_fd_sc_hd__o21ai_1 _13310_ (.A1(_05995_),
    .A2(_05921_),
    .B1(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__xor2_1 _13311_ (.A(_06044_),
    .B(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__nand2_1 _13312_ (.A(_06022_),
    .B(_06038_),
    .Y(_06049_));
 sky130_fd_sc_hd__o21ai_1 _13313_ (.A1(_06039_),
    .A2(_06048_),
    .B1(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__xnor2_1 _13314_ (.A(_06021_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__or2_1 _13315_ (.A(_05973_),
    .B(_05961_),
    .X(_06052_));
 sky130_fd_sc_hd__or3b_4 _13316_ (.A(_05939_),
    .B(_06052_),
    .C_N(_05922_),
    .X(_06053_));
 sky130_fd_sc_hd__nor2_1 _13317_ (.A(_05939_),
    .B(_05961_),
    .Y(_06054_));
 sky130_fd_sc_hd__inv_2 _13318_ (.A(_05973_),
    .Y(_06055_));
 sky130_fd_sc_hd__a21o_1 _13319_ (.A1(_05922_),
    .A2(_06054_),
    .B1(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__clkbuf_4 _13320_ (.A(_05947_),
    .X(_06057_));
 sky130_fd_sc_hd__a21o_1 _13321_ (.A1(_06053_),
    .A2(_06056_),
    .B1(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _13322_ (.A(_05923_),
    .B(_06054_),
    .Y(_06059_));
 sky130_fd_sc_hd__a21bo_1 _13323_ (.A1(_05923_),
    .A2(_05989_),
    .B1_N(_05983_),
    .X(_06060_));
 sky130_fd_sc_hd__clkbuf_4 _13324_ (.A(_05944_),
    .X(_06061_));
 sky130_fd_sc_hd__a21oi_2 _13325_ (.A1(_06059_),
    .A2(_06060_),
    .B1(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__inv_2 _13326_ (.A(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_1 _13327_ (.A(_06058_),
    .B(_06062_),
    .Y(_06064_));
 sky130_fd_sc_hd__nand2_4 _13328_ (.A(_05852_),
    .B(_05853_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_1 _13329_ (.A(_05752_),
    .B(_06053_),
    .Y(_06066_));
 sky130_fd_sc_hd__clkbuf_4 _13330_ (.A(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__nor2_1 _13331_ (.A(_06065_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__a2bb2o_1 _13332_ (.A1_N(_06058_),
    .A2_N(_06063_),
    .B1(_06064_),
    .B2(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__nor2_1 _13333_ (.A(_06057_),
    .B(_06067_),
    .Y(_06070_));
 sky130_fd_sc_hd__a21o_1 _13334_ (.A1(_06053_),
    .A2(_06056_),
    .B1(_06061_),
    .X(_06071_));
 sky130_fd_sc_hd__a21oi_1 _13335_ (.A1(_06059_),
    .A2(_06060_),
    .B1(_06045_),
    .Y(_06072_));
 sky130_fd_sc_hd__xnor2_1 _13336_ (.A(_06071_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__xor2_2 _13337_ (.A(_06070_),
    .B(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__nand2_1 _13338_ (.A(_06069_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__and2b_1 _13339_ (.A_N(_06044_),
    .B(_06047_),
    .X(_06076_));
 sky130_fd_sc_hd__a21oi_1 _13340_ (.A1(_06040_),
    .A2(_06043_),
    .B1(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__clkbuf_4 _13341_ (.A(_06045_),
    .X(_06078_));
 sky130_fd_sc_hd__and2_1 _13342_ (.A(_06053_),
    .B(_06056_),
    .X(_06079_));
 sky130_fd_sc_hd__clkbuf_4 _13343_ (.A(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__or2_1 _13344_ (.A(_06078_),
    .B(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__a2bb2o_1 _13345_ (.A1_N(_06063_),
    .A2_N(_06081_),
    .B1(_06073_),
    .B2(_06070_),
    .X(_06082_));
 sky130_fd_sc_hd__or2_1 _13346_ (.A(_06061_),
    .B(_06067_),
    .X(_06083_));
 sky130_fd_sc_hd__and2_1 _13347_ (.A(_06059_),
    .B(_06060_),
    .X(_06084_));
 sky130_fd_sc_hd__nor2_1 _13348_ (.A(_06041_),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__xnor2_1 _13349_ (.A(_06081_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__xnor2_1 _13350_ (.A(_06083_),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__xor2_1 _13351_ (.A(_06082_),
    .B(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__xnor2_1 _13352_ (.A(_06077_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__xnor2_1 _13353_ (.A(_06075_),
    .B(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__xnor2_1 _13354_ (.A(_06051_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__a21bo_1 _13355_ (.A1(_06036_),
    .A2(_06035_),
    .B1_N(_06030_),
    .X(_06092_));
 sky130_fd_sc_hd__a21oi_1 _13356_ (.A1(_05945_),
    .A2(_05949_),
    .B1(_05939_),
    .Y(_06093_));
 sky130_fd_sc_hd__o21bai_1 _13357_ (.A1(_05991_),
    .A2(_05975_),
    .B1_N(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__or3b_1 _13358_ (.A(_05920_),
    .B(_05975_),
    .C_N(_06093_),
    .X(_06095_));
 sky130_fd_sc_hd__a21oi_1 _13359_ (.A1(_05941_),
    .A2(_05980_),
    .B1(_05990_),
    .Y(_06096_));
 sky130_fd_sc_hd__nand3_1 _13360_ (.A(_06094_),
    .B(_06095_),
    .C(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__a21o_1 _13361_ (.A1(_06094_),
    .A2(_06095_),
    .B1(_06096_),
    .X(_06098_));
 sky130_fd_sc_hd__xnor2_1 _13362_ (.A(_06025_),
    .B(_06027_),
    .Y(_06099_));
 sky130_fd_sc_hd__or2_1 _13363_ (.A(_05823_),
    .B(_05973_),
    .X(_06100_));
 sky130_fd_sc_hd__or3_1 _13364_ (.A(_05946_),
    .B(_05961_),
    .C(_06007_),
    .X(_06101_));
 sky130_fd_sc_hd__or2_1 _13365_ (.A(_06100_),
    .B(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__nor2_1 _13366_ (.A(_05939_),
    .B(_06016_),
    .Y(_06103_));
 sky130_fd_sc_hd__xor2_1 _13367_ (.A(_06100_),
    .B(_06101_),
    .X(_06104_));
 sky130_fd_sc_hd__nand2_1 _13368_ (.A(_06103_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__nand3_1 _13369_ (.A(_06099_),
    .B(_06102_),
    .C(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__a21oi_1 _13370_ (.A1(_06102_),
    .A2(_06105_),
    .B1(_06099_),
    .Y(_06107_));
 sky130_fd_sc_hd__a31o_1 _13371_ (.A1(_06097_),
    .A2(_06098_),
    .A3(_06106_),
    .B1(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__and3_1 _13372_ (.A(_06037_),
    .B(_06092_),
    .C(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__a21oi_1 _13373_ (.A1(_06037_),
    .A2(_06092_),
    .B1(_06108_),
    .Y(_06110_));
 sky130_fd_sc_hd__nor2_1 _13374_ (.A(_06109_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__nor2_1 _13375_ (.A(_06061_),
    .B(_05940_),
    .Y(_06112_));
 sky130_fd_sc_hd__a21o_1 _13376_ (.A1(_05889_),
    .A2(_05900_),
    .B1(_05910_),
    .X(_06113_));
 sky130_fd_sc_hd__a21o_1 _13377_ (.A1(_05995_),
    .A2(_06113_),
    .B1(_05846_),
    .X(_06114_));
 sky130_fd_sc_hd__inv_2 _13378_ (.A(_06045_),
    .Y(_06115_));
 sky130_fd_sc_hd__or4b_2 _13379_ (.A(_05979_),
    .B(_05909_),
    .C(_05920_),
    .D_N(_05900_),
    .X(_06116_));
 sky130_fd_sc_hd__and3_1 _13380_ (.A(_06115_),
    .B(_05923_),
    .C(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__xnor2_2 _13381_ (.A(_06114_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__nand2_1 _13382_ (.A(_05923_),
    .B(_06116_),
    .Y(_06119_));
 sky130_fd_sc_hd__or3_1 _13383_ (.A(_06045_),
    .B(_06114_),
    .C(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__a21bo_1 _13384_ (.A1(_06112_),
    .A2(_06118_),
    .B1_N(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__a21boi_1 _13385_ (.A1(_06094_),
    .A2(_06096_),
    .B1_N(_06095_),
    .Y(_06122_));
 sky130_fd_sc_hd__o22ai_1 _13386_ (.A1(_06041_),
    .A2(_05991_),
    .B1(_05940_),
    .B2(_06078_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand3b_1 _13387_ (.A_N(_06122_),
    .B(_06046_),
    .C(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__a21bo_1 _13388_ (.A1(_06046_),
    .A2(_06123_),
    .B1_N(_06122_),
    .X(_06125_));
 sky130_fd_sc_hd__and3_1 _13389_ (.A(_06121_),
    .B(_06124_),
    .C(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__a21oi_1 _13390_ (.A1(_06124_),
    .A2(_06125_),
    .B1(_06121_),
    .Y(_06127_));
 sky130_fd_sc_hd__nor2_1 _13391_ (.A(_06126_),
    .B(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__a21o_1 _13392_ (.A1(_06111_),
    .A2(_06128_),
    .B1(_06109_),
    .X(_06129_));
 sky130_fd_sc_hd__xnor2_1 _13393_ (.A(_06039_),
    .B(_06048_),
    .Y(_06130_));
 sky130_fd_sc_hd__xnor2_1 _13394_ (.A(_06129_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__or2_1 _13395_ (.A(_05824_),
    .B(_06066_),
    .X(_06132_));
 sky130_fd_sc_hd__o22a_1 _13396_ (.A1(_06065_),
    .A2(_06080_),
    .B1(_06084_),
    .B2(_06057_),
    .X(_06133_));
 sky130_fd_sc_hd__clkbuf_4 _13397_ (.A(_06084_),
    .X(_06134_));
 sky130_fd_sc_hd__nor3_1 _13398_ (.A(_06065_),
    .B(_06058_),
    .C(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__o21ba_1 _13399_ (.A1(_06132_),
    .A2(_06133_),
    .B1_N(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__xor2_1 _13400_ (.A(_06068_),
    .B(_06064_),
    .X(_06137_));
 sky130_fd_sc_hd__or2b_1 _13401_ (.A(_06136_),
    .B_N(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__a21bo_1 _13402_ (.A1(_06121_),
    .A2(_06125_),
    .B1_N(_06124_),
    .X(_06139_));
 sky130_fd_sc_hd__xor2_1 _13403_ (.A(_06069_),
    .B(_06074_),
    .X(_06140_));
 sky130_fd_sc_hd__xnor2_1 _13404_ (.A(_06139_),
    .B(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__xor2_1 _13405_ (.A(_06138_),
    .B(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__and2b_1 _13406_ (.A_N(_06130_),
    .B(_06129_),
    .X(_06143_));
 sky130_fd_sc_hd__a21o_1 _13407_ (.A1(_06131_),
    .A2(_06142_),
    .B1(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__and2b_1 _13408_ (.A_N(_06091_),
    .B(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(_06139_),
    .B(_06140_),
    .Y(_06146_));
 sky130_fd_sc_hd__o21a_1 _13410_ (.A1(_06138_),
    .A2(_06141_),
    .B1(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__xnor2_1 _13411_ (.A(_06144_),
    .B(_06091_),
    .Y(_06148_));
 sky130_fd_sc_hd__and2b_1 _13412_ (.A_N(_06147_),
    .B(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__nor2_1 _13413_ (.A(_06145_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__and2b_1 _13414_ (.A_N(_06021_),
    .B(_06050_),
    .X(_06151_));
 sky130_fd_sc_hd__a21oi_1 _13415_ (.A1(_06051_),
    .A2(_06090_),
    .B1(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_4 _13416_ (.A(_05988_),
    .B(_05980_),
    .Y(_06153_));
 sky130_fd_sc_hd__and3_1 _13417_ (.A(_05752_),
    .B(_06153_),
    .C(_05976_),
    .X(_06154_));
 sky130_fd_sc_hd__o22a_1 _13418_ (.A1(_06015_),
    .A2(_06031_),
    .B1(_05982_),
    .B2(_05974_),
    .X(_06155_));
 sky130_fd_sc_hd__or2_1 _13419_ (.A(_06154_),
    .B(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__nor2_1 _13420_ (.A(_05978_),
    .B(_05942_),
    .Y(_06157_));
 sky130_fd_sc_hd__a21bo_1 _13421_ (.A1(_06002_),
    .A2(_05976_),
    .B1_N(_06004_),
    .X(_06158_));
 sky130_fd_sc_hd__and2_1 _13422_ (.A(_05995_),
    .B(_06113_),
    .X(_06159_));
 sky130_fd_sc_hd__nor2_1 _13423_ (.A(_05983_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__clkbuf_4 _13424_ (.A(_06119_),
    .X(_06161_));
 sky130_fd_sc_hd__nor2_1 _13425_ (.A(_05978_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__xor2_1 _13426_ (.A(_06160_),
    .B(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__nor2_1 _13427_ (.A(_05991_),
    .B(_05978_),
    .Y(_06164_));
 sky130_fd_sc_hd__xnor2_1 _13428_ (.A(_06163_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__xnor2_1 _13429_ (.A(_06158_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__xnor2_1 _13430_ (.A(_06157_),
    .B(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__nor2_1 _13431_ (.A(_06156_),
    .B(_06167_),
    .Y(_06168_));
 sky130_fd_sc_hd__and2_1 _13432_ (.A(_06156_),
    .B(_06167_),
    .X(_06169_));
 sky130_fd_sc_hd__or2_1 _13433_ (.A(_06168_),
    .B(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__a32o_1 _13434_ (.A1(_06004_),
    .A2(_06005_),
    .A3(_06019_),
    .B1(_06020_),
    .B2(_06001_),
    .X(_06171_));
 sky130_fd_sc_hd__xor2_1 _13435_ (.A(_06170_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__nand2_1 _13436_ (.A(_06082_),
    .B(_06087_),
    .Y(_06173_));
 sky130_fd_sc_hd__and2b_1 _13437_ (.A_N(_05943_),
    .B(_06000_),
    .X(_06174_));
 sky130_fd_sc_hd__or2_1 _13438_ (.A(_05998_),
    .B(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__clkinv_2 _13439_ (.A(_06080_),
    .Y(_06176_));
 sky130_fd_sc_hd__and3_1 _13440_ (.A(_06115_),
    .B(_06176_),
    .C(_06085_),
    .X(_06177_));
 sky130_fd_sc_hd__and2b_1 _13441_ (.A_N(_06083_),
    .B(_06086_),
    .X(_06178_));
 sky130_fd_sc_hd__or2_1 _13442_ (.A(_06078_),
    .B(_06067_),
    .X(_06179_));
 sky130_fd_sc_hd__o22a_1 _13443_ (.A1(_06041_),
    .A2(_06080_),
    .B1(_06084_),
    .B2(_05990_),
    .X(_06180_));
 sky130_fd_sc_hd__a31oi_1 _13444_ (.A1(_05910_),
    .A2(_06176_),
    .A3(_06085_),
    .B1(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__xnor2_1 _13445_ (.A(_06179_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__o21ai_1 _13446_ (.A1(_06177_),
    .A2(_06178_),
    .B1(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__or3_1 _13447_ (.A(_06177_),
    .B(_06178_),
    .C(_06182_),
    .X(_06184_));
 sky130_fd_sc_hd__and2_1 _13448_ (.A(_06183_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__xnor2_1 _13449_ (.A(_06175_),
    .B(_06185_),
    .Y(_06186_));
 sky130_fd_sc_hd__xor2_1 _13450_ (.A(_06173_),
    .B(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__xnor2_1 _13451_ (.A(_06172_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__xnor2_1 _13452_ (.A(_06152_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__and2b_1 _13453_ (.A_N(_06077_),
    .B(_06088_),
    .X(_06190_));
 sky130_fd_sc_hd__a31oi_2 _13454_ (.A1(_06069_),
    .A2(_06074_),
    .A3(_06089_),
    .B1(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__xnor2_1 _13455_ (.A(_06189_),
    .B(_06191_),
    .Y(_06192_));
 sky130_fd_sc_hd__and2b_1 _13456_ (.A_N(_06150_),
    .B(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__or2b_1 _13457_ (.A(_06152_),
    .B_N(_06188_),
    .X(_06194_));
 sky130_fd_sc_hd__or2b_1 _13458_ (.A(_06191_),
    .B_N(_06189_),
    .X(_06195_));
 sky130_fd_sc_hd__nand2_1 _13459_ (.A(_06194_),
    .B(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__and2b_1 _13460_ (.A_N(_06170_),
    .B(_06171_),
    .X(_06197_));
 sky130_fd_sc_hd__and2b_1 _13461_ (.A_N(_06172_),
    .B(_06187_),
    .X(_06198_));
 sky130_fd_sc_hd__nand2_1 _13462_ (.A(_05752_),
    .B(_06153_),
    .Y(_06199_));
 sky130_fd_sc_hd__a22o_1 _13463_ (.A1(_06160_),
    .A2(_06162_),
    .B1(_06163_),
    .B2(_06164_),
    .X(_06200_));
 sky130_fd_sc_hd__nand2_2 _13464_ (.A(_05923_),
    .B(_05989_),
    .Y(_06201_));
 sky130_fd_sc_hd__nor2_1 _13465_ (.A(_05974_),
    .B(_06161_),
    .Y(_06202_));
 sky130_fd_sc_hd__o22a_1 _13466_ (.A1(_05974_),
    .A2(_06159_),
    .B1(_06161_),
    .B2(_05983_),
    .X(_06203_));
 sky130_fd_sc_hd__a21o_1 _13467_ (.A1(_06160_),
    .A2(_06202_),
    .B1(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__xor2_1 _13468_ (.A(_06201_),
    .B(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__xnor2_1 _13469_ (.A(_06154_),
    .B(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__xnor2_1 _13470_ (.A(_06200_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__xnor2_1 _13471_ (.A(_06199_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__xnor2_1 _13472_ (.A(_06168_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__or2b_1 _13473_ (.A(_06165_),
    .B_N(_06158_),
    .X(_06210_));
 sky130_fd_sc_hd__a21bo_1 _13474_ (.A1(_06157_),
    .A2(_06166_),
    .B1_N(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__and3_1 _13475_ (.A(_05910_),
    .B(_06176_),
    .C(_06085_),
    .X(_06212_));
 sky130_fd_sc_hd__and2b_1 _13476_ (.A_N(_06179_),
    .B(_06181_),
    .X(_06213_));
 sky130_fd_sc_hd__or2_1 _13477_ (.A(_06041_),
    .B(_06067_),
    .X(_06214_));
 sky130_fd_sc_hd__nor2_1 _13478_ (.A(_05990_),
    .B(_06134_),
    .Y(_06215_));
 sky130_fd_sc_hd__o22a_1 _13479_ (.A1(_05990_),
    .A2(_06080_),
    .B1(_06084_),
    .B2(_05991_),
    .X(_06216_));
 sky130_fd_sc_hd__a31oi_1 _13480_ (.A1(_05921_),
    .A2(_06176_),
    .A3(_06215_),
    .B1(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__xnor2_1 _13481_ (.A(_06214_),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__o21ai_2 _13482_ (.A1(_06212_),
    .A2(_06213_),
    .B1(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__or3_1 _13483_ (.A(_06212_),
    .B(_06213_),
    .C(_06218_),
    .X(_06220_));
 sky130_fd_sc_hd__and2_1 _13484_ (.A(_06219_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__xnor2_1 _13485_ (.A(_06211_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__xor2_1 _13486_ (.A(_06183_),
    .B(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__xnor2_1 _13487_ (.A(_06209_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__o21ai_1 _13488_ (.A1(_06197_),
    .A2(_06198_),
    .B1(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__or3_1 _13489_ (.A(_06197_),
    .B(_06198_),
    .C(_06224_),
    .X(_06226_));
 sky130_fd_sc_hd__and2_1 _13490_ (.A(_06225_),
    .B(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__nor2_1 _13491_ (.A(_06173_),
    .B(_06186_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21oi_1 _13492_ (.A1(_06175_),
    .A2(_06185_),
    .B1(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__xor2_1 _13493_ (.A(_06227_),
    .B(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__xnor2_1 _13494_ (.A(_06196_),
    .B(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__and2b_1 _13495_ (.A_N(_06230_),
    .B(_06196_),
    .X(_06232_));
 sky130_fd_sc_hd__or2b_1 _13496_ (.A(_06229_),
    .B_N(_06227_),
    .X(_06233_));
 sky130_fd_sc_hd__and2b_1 _13497_ (.A_N(_06209_),
    .B(_06223_),
    .X(_06234_));
 sky130_fd_sc_hd__a21o_1 _13498_ (.A1(_06168_),
    .A2(_06208_),
    .B1(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__and3_1 _13499_ (.A(_05752_),
    .B(_06153_),
    .C(_06207_),
    .X(_06236_));
 sky130_fd_sc_hd__nand2_1 _13500_ (.A(_06160_),
    .B(_06202_),
    .Y(_06237_));
 sky130_fd_sc_hd__or2_1 _13501_ (.A(_06201_),
    .B(_06204_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_4 _13502_ (.A(_06015_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_4 _13503_ (.A(_06159_),
    .X(_06240_));
 sky130_fd_sc_hd__o21bai_1 _13504_ (.A1(_06239_),
    .A2(_06240_),
    .B1_N(_06202_),
    .Y(_06241_));
 sky130_fd_sc_hd__or3_1 _13505_ (.A(_05974_),
    .B(_06240_),
    .C(_06161_),
    .X(_06242_));
 sky130_fd_sc_hd__nand2_1 _13506_ (.A(_06241_),
    .B(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__or3_1 _13507_ (.A(_05983_),
    .B(_05940_),
    .C(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_4 _13508_ (.A(_05940_),
    .X(_06245_));
 sky130_fd_sc_hd__o21ai_1 _13509_ (.A1(_05983_),
    .A2(_06245_),
    .B1(_06243_),
    .Y(_06246_));
 sky130_fd_sc_hd__nand2_1 _13510_ (.A(_06244_),
    .B(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__a21oi_2 _13511_ (.A1(_06237_),
    .A2(_06238_),
    .B1(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__and3_1 _13512_ (.A(_06237_),
    .B(_06238_),
    .C(_06247_),
    .X(_06249_));
 sky130_fd_sc_hd__nor2_1 _13513_ (.A(_06248_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_1 _13514_ (.A(_06236_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__or2_1 _13515_ (.A(_06236_),
    .B(_06250_),
    .X(_06252_));
 sky130_fd_sc_hd__and2_1 _13516_ (.A(_06251_),
    .B(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__or2b_1 _13517_ (.A(_06206_),
    .B_N(_06200_),
    .X(_06254_));
 sky130_fd_sc_hd__a21bo_1 _13518_ (.A1(_06154_),
    .A2(_06205_),
    .B1_N(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__and3_1 _13519_ (.A(_05921_),
    .B(_06176_),
    .C(_06215_),
    .X(_06256_));
 sky130_fd_sc_hd__and2b_1 _13520_ (.A_N(_06214_),
    .B(_06217_),
    .X(_06257_));
 sky130_fd_sc_hd__or2_1 _13521_ (.A(_05990_),
    .B(_06067_),
    .X(_06258_));
 sky130_fd_sc_hd__and4bb_1 _13522_ (.A_N(_06080_),
    .B_N(_06134_),
    .C(_05921_),
    .D(_05989_),
    .X(_06259_));
 sky130_fd_sc_hd__o22a_1 _13523_ (.A1(_05991_),
    .A2(_06080_),
    .B1(_06134_),
    .B2(_05978_),
    .X(_06260_));
 sky130_fd_sc_hd__nor2_1 _13524_ (.A(_06259_),
    .B(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__xnor2_1 _13525_ (.A(_06258_),
    .B(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__o21ai_1 _13526_ (.A1(_06256_),
    .A2(_06257_),
    .B1(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__or3_1 _13527_ (.A(_06256_),
    .B(_06257_),
    .C(_06262_),
    .X(_06264_));
 sky130_fd_sc_hd__and2_1 _13528_ (.A(_06263_),
    .B(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__xnor2_1 _13529_ (.A(_06255_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__xor2_1 _13530_ (.A(_06219_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__xnor2_1 _13531_ (.A(_06253_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__xnor2_1 _13532_ (.A(_06235_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__nor2_1 _13533_ (.A(_06183_),
    .B(_06222_),
    .Y(_06270_));
 sky130_fd_sc_hd__a21oi_1 _13534_ (.A1(_06211_),
    .A2(_06221_),
    .B1(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__xor2_1 _13535_ (.A(_06269_),
    .B(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__a21oi_1 _13536_ (.A1(_06225_),
    .A2(_06233_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__and3_1 _13537_ (.A(_06225_),
    .B(_06233_),
    .C(_06272_),
    .X(_06274_));
 sky130_fd_sc_hd__nor2_1 _13538_ (.A(_06273_),
    .B(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__xor2_1 _13539_ (.A(_06232_),
    .B(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__and3_1 _13540_ (.A(_06193_),
    .B(_06231_),
    .C(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__xor2_1 _13541_ (.A(_06193_),
    .B(_06231_),
    .X(_06278_));
 sky130_fd_sc_hd__xnor2_2 _13542_ (.A(_06150_),
    .B(_06192_),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_1 _13543_ (.A(_06135_),
    .B(_06133_),
    .Y(_06280_));
 sky130_fd_sc_hd__xor2_2 _13544_ (.A(_06132_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__or2_1 _13545_ (.A(_06065_),
    .B(_06134_),
    .X(_06282_));
 sky130_fd_sc_hd__or3_2 _13546_ (.A(_05824_),
    .B(_06080_),
    .C(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__xor2_1 _13547_ (.A(_06136_),
    .B(_06137_),
    .X(_06284_));
 sky130_fd_sc_hd__a21oi_1 _13548_ (.A1(_05945_),
    .A2(_05949_),
    .B1(_05990_),
    .Y(_06285_));
 sky130_fd_sc_hd__and3b_1 _13549_ (.A_N(_05975_),
    .B(_06285_),
    .C(_05921_),
    .X(_06286_));
 sky130_fd_sc_hd__o22a_1 _13550_ (.A1(_05990_),
    .A2(_05975_),
    .B1(_05984_),
    .B2(_05991_),
    .X(_06287_));
 sky130_fd_sc_hd__nor3_1 _13551_ (.A(_05988_),
    .B(_06287_),
    .C(_06286_),
    .Y(_06288_));
 sky130_fd_sc_hd__or2_1 _13552_ (.A(_06286_),
    .B(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__xor2_2 _13553_ (.A(_06112_),
    .B(_06118_),
    .X(_06290_));
 sky130_fd_sc_hd__xnor2_2 _13554_ (.A(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__a21o_1 _13555_ (.A1(_05995_),
    .A2(_06113_),
    .B1(_06061_),
    .X(_06292_));
 sky130_fd_sc_hd__nor2_1 _13556_ (.A(_06057_),
    .B(_05940_),
    .Y(_06293_));
 sky130_fd_sc_hd__a21o_1 _13557_ (.A1(_05995_),
    .A2(_06113_),
    .B1(_06045_),
    .X(_06294_));
 sky130_fd_sc_hd__and3_1 _13558_ (.A(_05888_),
    .B(_05923_),
    .C(_06116_),
    .X(_06295_));
 sky130_fd_sc_hd__xnor2_1 _13559_ (.A(_06294_),
    .B(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(_06293_),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__o31a_1 _13561_ (.A1(_06078_),
    .A2(_06161_),
    .A3(_06292_),
    .B1(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__nand2_1 _13562_ (.A(_06289_),
    .B(_06290_),
    .Y(_06299_));
 sky130_fd_sc_hd__o21a_1 _13563_ (.A1(_06291_),
    .A2(_06298_),
    .B1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__xnor2_1 _13564_ (.A(_06284_),
    .B(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__o32a_1 _13565_ (.A1(_06281_),
    .A2(_06283_),
    .A3(_06301_),
    .B1(_06300_),
    .B2(_06284_),
    .X(_06302_));
 sky130_fd_sc_hd__xnor2_1 _13566_ (.A(_06131_),
    .B(_06142_),
    .Y(_06303_));
 sky130_fd_sc_hd__xnor2_2 _13567_ (.A(_06111_),
    .B(_06128_),
    .Y(_06304_));
 sky130_fd_sc_hd__xor2_2 _13568_ (.A(_06291_),
    .B(_06298_),
    .X(_06305_));
 sky130_fd_sc_hd__and2_1 _13569_ (.A(_06097_),
    .B(_06098_),
    .X(_06306_));
 sky130_fd_sc_hd__and2b_1 _13570_ (.A_N(_06107_),
    .B(_06106_),
    .X(_06307_));
 sky130_fd_sc_hd__xnor2_2 _13571_ (.A(_06306_),
    .B(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__xnor2_1 _13572_ (.A(_06103_),
    .B(_06104_),
    .Y(_06309_));
 sky130_fd_sc_hd__or2_1 _13573_ (.A(_05823_),
    .B(_05939_),
    .X(_06310_));
 sky130_fd_sc_hd__or2_1 _13574_ (.A(_05920_),
    .B(_06016_),
    .X(_06311_));
 sky130_fd_sc_hd__or2_1 _13575_ (.A(_05823_),
    .B(_05961_),
    .X(_06312_));
 sky130_fd_sc_hd__or3_2 _13576_ (.A(_05946_),
    .B(_05939_),
    .C(_06007_),
    .X(_06313_));
 sky130_fd_sc_hd__xnor2_1 _13577_ (.A(_06312_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__o22a_1 _13578_ (.A1(_06101_),
    .A2(_06310_),
    .B1(_06311_),
    .B2(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__nand2_1 _13579_ (.A(_06309_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__o21a_1 _13580_ (.A1(_06287_),
    .A2(_06286_),
    .B1(_05988_),
    .X(_06317_));
 sky130_fd_sc_hd__nor2_1 _13581_ (.A(_06288_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__nor2_1 _13582_ (.A(_06309_),
    .B(_06315_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21o_1 _13583_ (.A1(_06316_),
    .A2(_06318_),
    .B1(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__xnor2_2 _13584_ (.A(_06308_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__and2b_1 _13585_ (.A_N(_06308_),
    .B(_06320_),
    .X(_06322_));
 sky130_fd_sc_hd__a21oi_1 _13586_ (.A1(_06305_),
    .A2(_06321_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2_1 _13587_ (.A(_06304_),
    .B(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__nor2_1 _13588_ (.A(_06281_),
    .B(_06283_),
    .Y(_06325_));
 sky130_fd_sc_hd__xnor2_1 _13589_ (.A(_06325_),
    .B(_06301_),
    .Y(_06326_));
 sky130_fd_sc_hd__nor2_1 _13590_ (.A(_06304_),
    .B(_06323_),
    .Y(_06327_));
 sky130_fd_sc_hd__a21oi_1 _13591_ (.A1(_06324_),
    .A2(_06326_),
    .B1(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__xnor2_1 _13592_ (.A(_06303_),
    .B(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__nor2_1 _13593_ (.A(_06303_),
    .B(_06328_),
    .Y(_06330_));
 sky130_fd_sc_hd__o21ba_1 _13594_ (.A1(_06302_),
    .A2(_06329_),
    .B1_N(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__xnor2_1 _13595_ (.A(_06148_),
    .B(_06147_),
    .Y(_06332_));
 sky130_fd_sc_hd__and2b_1 _13596_ (.A_N(_06331_),
    .B(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__and2_1 _13597_ (.A(_06279_),
    .B(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__nand2_1 _13598_ (.A(_06278_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_1 _13599_ (.A(_06302_),
    .B(_06329_),
    .Y(_06336_));
 sky130_fd_sc_hd__xnor2_1 _13600_ (.A(_06293_),
    .B(_06296_),
    .Y(_06337_));
 sky130_fd_sc_hd__xnor2_1 _13601_ (.A(_05988_),
    .B(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__a21oi_2 _13602_ (.A1(_05995_),
    .A2(_06113_),
    .B1(_06057_),
    .Y(_06339_));
 sky130_fd_sc_hd__nor2_1 _13603_ (.A(_06065_),
    .B(_05940_),
    .Y(_06340_));
 sky130_fd_sc_hd__and3_1 _13604_ (.A(_05877_),
    .B(_05923_),
    .C(_06116_),
    .X(_06341_));
 sky130_fd_sc_hd__xnor2_1 _13605_ (.A(_06292_),
    .B(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__a22o_1 _13606_ (.A1(_06295_),
    .A2(_06339_),
    .B1(_06340_),
    .B2(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__and2b_1 _13607_ (.A_N(_06338_),
    .B(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__o21ba_1 _13608_ (.A1(_05988_),
    .A2(_06337_),
    .B1_N(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__xnor2_1 _13609_ (.A(_06281_),
    .B(_06283_),
    .Y(_06346_));
 sky130_fd_sc_hd__nor2_1 _13610_ (.A(_06345_),
    .B(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__xnor2_1 _13611_ (.A(_06304_),
    .B(_06323_),
    .Y(_06348_));
 sky130_fd_sc_hd__xnor2_1 _13612_ (.A(_06348_),
    .B(_06326_),
    .Y(_06349_));
 sky130_fd_sc_hd__xnor2_1 _13613_ (.A(_06345_),
    .B(_06346_),
    .Y(_06350_));
 sky130_fd_sc_hd__xor2_2 _13614_ (.A(_06305_),
    .B(_06321_),
    .X(_06351_));
 sky130_fd_sc_hd__xnor2_1 _13615_ (.A(_06338_),
    .B(_06343_),
    .Y(_06352_));
 sky130_fd_sc_hd__or2b_1 _13616_ (.A(_06319_),
    .B_N(_06316_),
    .X(_06353_));
 sky130_fd_sc_hd__xnor2_1 _13617_ (.A(_06353_),
    .B(_06318_),
    .Y(_06354_));
 sky130_fd_sc_hd__xnor2_1 _13618_ (.A(_06311_),
    .B(_06314_),
    .Y(_06355_));
 sky130_fd_sc_hd__or2_2 _13619_ (.A(_05823_),
    .B(_05920_),
    .X(_06356_));
 sky130_fd_sc_hd__or2_1 _13620_ (.A(_05990_),
    .B(_06016_),
    .X(_06357_));
 sky130_fd_sc_hd__o21a_1 _13621_ (.A1(_05920_),
    .A2(_06009_),
    .B1(_06310_),
    .X(_06358_));
 sky130_fd_sc_hd__o22a_1 _13622_ (.A1(_06313_),
    .A2(_06356_),
    .B1(_06357_),
    .B2(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__xor2_1 _13623_ (.A(_06355_),
    .B(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__or3_1 _13624_ (.A(_05846_),
    .B(_05975_),
    .C(_06285_),
    .X(_06361_));
 sky130_fd_sc_hd__o21ai_1 _13625_ (.A1(_06041_),
    .A2(_06031_),
    .B1(_06285_),
    .Y(_06362_));
 sky130_fd_sc_hd__a211o_1 _13626_ (.A1(_06361_),
    .A2(_06362_),
    .B1(_06078_),
    .C1(_05982_),
    .X(_06363_));
 sky130_fd_sc_hd__o211ai_1 _13627_ (.A1(_06078_),
    .A2(_05982_),
    .B1(_06361_),
    .C1(_06362_),
    .Y(_06364_));
 sky130_fd_sc_hd__and3_1 _13628_ (.A(_06360_),
    .B(_06363_),
    .C(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__o21ba_1 _13629_ (.A1(_06355_),
    .A2(_06359_),
    .B1_N(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__xnor2_1 _13630_ (.A(_06354_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__and2b_1 _13631_ (.A_N(_06366_),
    .B(_06354_),
    .X(_06368_));
 sky130_fd_sc_hd__a21o_1 _13632_ (.A1(_06352_),
    .A2(_06367_),
    .B1(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__nor2_1 _13633_ (.A(_06351_),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nand2_1 _13634_ (.A(_06351_),
    .B(_06369_),
    .Y(_06371_));
 sky130_fd_sc_hd__o21a_1 _13635_ (.A1(_06350_),
    .A2(_06370_),
    .B1(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__xnor2_2 _13636_ (.A(_06349_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__or2b_1 _13637_ (.A(_06372_),
    .B_N(_06349_),
    .X(_06374_));
 sky130_fd_sc_hd__a21boi_2 _13638_ (.A1(_06347_),
    .A2(_06373_),
    .B1_N(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__xor2_1 _13639_ (.A(_06332_),
    .B(_06331_),
    .X(_06376_));
 sky130_fd_sc_hd__nor3_1 _13640_ (.A(_06336_),
    .B(_06375_),
    .C(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_1 _13641_ (.A(_06279_),
    .B(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__xnor2_2 _13642_ (.A(_06347_),
    .B(_06373_),
    .Y(_06379_));
 sky130_fd_sc_hd__xnor2_1 _13643_ (.A(_06340_),
    .B(_06342_),
    .Y(_06380_));
 sky130_fd_sc_hd__xnor2_1 _13644_ (.A(_05988_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__inv_2 _13645_ (.A(_06065_),
    .Y(_06382_));
 sky130_fd_sc_hd__and3_1 _13646_ (.A(_06382_),
    .B(_05923_),
    .C(_06116_),
    .X(_06383_));
 sky130_fd_sc_hd__or2_1 _13647_ (.A(_05824_),
    .B(_05940_),
    .X(_06384_));
 sky130_fd_sc_hd__xnor2_1 _13648_ (.A(_06339_),
    .B(_06383_),
    .Y(_06385_));
 sky130_fd_sc_hd__o2bb2ai_1 _13649_ (.A1_N(_06339_),
    .A2_N(_06383_),
    .B1(_06384_),
    .B2(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__and2b_1 _13650_ (.A_N(_06381_),
    .B(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__o21bai_1 _13651_ (.A1(_05988_),
    .A2(_06380_),
    .B1_N(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__o21ai_1 _13652_ (.A1(_05824_),
    .A2(_06080_),
    .B1(_06282_),
    .Y(_06389_));
 sky130_fd_sc_hd__and2_1 _13653_ (.A(_06283_),
    .B(_06389_),
    .X(_06390_));
 sky130_fd_sc_hd__and2_1 _13654_ (.A(_06388_),
    .B(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__xor2_1 _13655_ (.A(_06351_),
    .B(_06369_),
    .X(_06392_));
 sky130_fd_sc_hd__xnor2_1 _13656_ (.A(_06350_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__xnor2_1 _13657_ (.A(_06388_),
    .B(_06390_),
    .Y(_06394_));
 sky130_fd_sc_hd__xnor2_1 _13658_ (.A(_06352_),
    .B(_06367_),
    .Y(_06395_));
 sky130_fd_sc_hd__xnor2_1 _13659_ (.A(_06381_),
    .B(_06386_),
    .Y(_06396_));
 sky130_fd_sc_hd__a21oi_1 _13660_ (.A1(_06363_),
    .A2(_06364_),
    .B1(_06360_),
    .Y(_06397_));
 sky130_fd_sc_hd__or2_1 _13661_ (.A(_06365_),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__o21bai_1 _13662_ (.A1(_06313_),
    .A2(_06356_),
    .B1_N(_06358_),
    .Y(_06399_));
 sky130_fd_sc_hd__xnor2_1 _13663_ (.A(_06357_),
    .B(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__or2_1 _13664_ (.A(_05990_),
    .B(_06009_),
    .X(_06401_));
 sky130_fd_sc_hd__or2_1 _13665_ (.A(_06041_),
    .B(_06016_),
    .X(_06402_));
 sky130_fd_sc_hd__xnor2_1 _13666_ (.A(_06356_),
    .B(_06401_),
    .Y(_06403_));
 sky130_fd_sc_hd__o22a_1 _13667_ (.A1(_06356_),
    .A2(_06401_),
    .B1(_06402_),
    .B2(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__xnor2_1 _13668_ (.A(_06400_),
    .B(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _13669_ (.A(_05856_),
    .B(_05877_),
    .Y(_06406_));
 sky130_fd_sc_hd__or2_1 _13670_ (.A(_06406_),
    .B(_06078_),
    .X(_06407_));
 sky130_fd_sc_hd__nand2_1 _13671_ (.A(_06061_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__or2_1 _13672_ (.A(_06041_),
    .B(_06406_),
    .X(_06409_));
 sky130_fd_sc_hd__xor2_1 _13673_ (.A(_06408_),
    .B(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__nor2_1 _13674_ (.A(_06400_),
    .B(_06404_),
    .Y(_06411_));
 sky130_fd_sc_hd__o21ba_1 _13675_ (.A1(_06405_),
    .A2(_06410_),
    .B1_N(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__xor2_1 _13676_ (.A(_06398_),
    .B(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__nor2_1 _13677_ (.A(_06398_),
    .B(_06412_),
    .Y(_06414_));
 sky130_fd_sc_hd__a21oi_1 _13678_ (.A1(_06396_),
    .A2(_06413_),
    .B1(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__xnor2_1 _13679_ (.A(_06395_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__or2_1 _13680_ (.A(_06395_),
    .B(_06415_),
    .X(_06417_));
 sky130_fd_sc_hd__o21a_1 _13681_ (.A1(_06394_),
    .A2(_06416_),
    .B1(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__xnor2_1 _13682_ (.A(_06393_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__and2b_1 _13683_ (.A_N(_06418_),
    .B(_06393_),
    .X(_06420_));
 sky130_fd_sc_hd__a21oi_2 _13684_ (.A1(_06391_),
    .A2(_06419_),
    .B1(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__nor2_1 _13685_ (.A(_06379_),
    .B(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__xor2_1 _13686_ (.A(_06336_),
    .B(_06375_),
    .X(_06423_));
 sky130_fd_sc_hd__and2_1 _13687_ (.A(_06422_),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__or2b_1 _13688_ (.A(_06376_),
    .B_N(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__xnor2_2 _13689_ (.A(_06379_),
    .B(_06421_),
    .Y(_06426_));
 sky130_fd_sc_hd__xnor2_1 _13690_ (.A(_06394_),
    .B(_06416_),
    .Y(_06427_));
 sky130_fd_sc_hd__or2_1 _13691_ (.A(_05824_),
    .B(_06134_),
    .X(_06428_));
 sky130_fd_sc_hd__xnor2_1 _13692_ (.A(_06384_),
    .B(_06385_),
    .Y(_06429_));
 sky130_fd_sc_hd__a21oi_1 _13693_ (.A1(_05945_),
    .A2(_06409_),
    .B1(_06078_),
    .Y(_06430_));
 sky130_fd_sc_hd__xor2_1 _13694_ (.A(_06429_),
    .B(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_1 _13695_ (.A(_05824_),
    .B(_06240_),
    .Y(_06432_));
 sky130_fd_sc_hd__nand2_1 _13696_ (.A(_06383_),
    .B(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__or2b_1 _13697_ (.A(_06429_),
    .B_N(_06430_),
    .X(_06434_));
 sky130_fd_sc_hd__o21a_1 _13698_ (.A1(_06431_),
    .A2(_06433_),
    .B1(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__or2_1 _13699_ (.A(_06428_),
    .B(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__nand2_1 _13700_ (.A(_06428_),
    .B(_06435_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand2_1 _13701_ (.A(_06436_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__xor2_1 _13702_ (.A(_06396_),
    .B(_06413_),
    .X(_06439_));
 sky130_fd_sc_hd__xor2_1 _13703_ (.A(_06431_),
    .B(_06433_),
    .X(_06440_));
 sky130_fd_sc_hd__xor2_1 _13704_ (.A(_06405_),
    .B(_06410_),
    .X(_06441_));
 sky130_fd_sc_hd__xnor2_1 _13705_ (.A(_06402_),
    .B(_06403_),
    .Y(_06442_));
 sky130_fd_sc_hd__or2_1 _13706_ (.A(_05823_),
    .B(_05909_),
    .X(_06443_));
 sky130_fd_sc_hd__or2_1 _13707_ (.A(_05846_),
    .B(_06009_),
    .X(_06444_));
 sky130_fd_sc_hd__xnor2_1 _13708_ (.A(_06443_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__or2_1 _13709_ (.A(_06443_),
    .B(_06444_),
    .X(_06446_));
 sky130_fd_sc_hd__o31a_1 _13710_ (.A1(_06078_),
    .A2(_06016_),
    .A3(_06445_),
    .B1(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__xor2_1 _13711_ (.A(_06442_),
    .B(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__nor2_1 _13712_ (.A(_06057_),
    .B(_05982_),
    .Y(_06449_));
 sky130_fd_sc_hd__mux2_1 _13713_ (.A0(_06041_),
    .A1(_06449_),
    .S(_06407_),
    .X(_06450_));
 sky130_fd_sc_hd__a2bb2o_1 _13714_ (.A1_N(_06442_),
    .A2_N(_06447_),
    .B1(_06448_),
    .B2(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__or2_1 _13715_ (.A(_06441_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__and2_1 _13716_ (.A(_06441_),
    .B(_06451_),
    .X(_06453_));
 sky130_fd_sc_hd__a21oi_1 _13717_ (.A1(_06440_),
    .A2(_06452_),
    .B1(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__xor2_1 _13718_ (.A(_06439_),
    .B(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__or2b_1 _13719_ (.A(_06454_),
    .B_N(_06439_),
    .X(_06456_));
 sky130_fd_sc_hd__o21ai_1 _13720_ (.A1(_06438_),
    .A2(_06455_),
    .B1(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__or2b_1 _13721_ (.A(_06427_),
    .B_N(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__xnor2_1 _13722_ (.A(_06427_),
    .B(_06457_),
    .Y(_06459_));
 sky130_fd_sc_hd__or2b_1 _13723_ (.A(_06436_),
    .B_N(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__xnor2_1 _13724_ (.A(_06391_),
    .B(_06419_),
    .Y(_06461_));
 sky130_fd_sc_hd__a21o_1 _13725_ (.A1(_06458_),
    .A2(_06460_),
    .B1(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__nor2_1 _13726_ (.A(_06426_),
    .B(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(_06423_),
    .B(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__xor2_1 _13728_ (.A(_06436_),
    .B(_06459_),
    .X(_06465_));
 sky130_fd_sc_hd__or2b_1 _13729_ (.A(_06453_),
    .B_N(_06452_),
    .X(_06466_));
 sky130_fd_sc_hd__xor2_1 _13730_ (.A(_06440_),
    .B(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__xor2_1 _13731_ (.A(_06448_),
    .B(_06450_),
    .X(_06468_));
 sky130_fd_sc_hd__or3_1 _13732_ (.A(_06057_),
    .B(_06045_),
    .C(_05945_),
    .X(_06469_));
 sky130_fd_sc_hd__o21ai_1 _13733_ (.A1(_06057_),
    .A2(_06031_),
    .B1(_05945_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand4_1 _13734_ (.A(_06382_),
    .B(_06153_),
    .C(_06469_),
    .D(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__a22o_1 _13735_ (.A1(_06382_),
    .A2(_06153_),
    .B1(_06469_),
    .B2(_06470_),
    .X(_06472_));
 sky130_fd_sc_hd__nor2_1 _13736_ (.A(_06045_),
    .B(_06016_),
    .Y(_06473_));
 sky130_fd_sc_hd__xnor2_1 _13737_ (.A(_06473_),
    .B(_06445_),
    .Y(_06474_));
 sky130_fd_sc_hd__nor2_1 _13738_ (.A(_05846_),
    .B(_05823_),
    .Y(_06475_));
 sky130_fd_sc_hd__nor2_1 _13739_ (.A(_06045_),
    .B(_06009_),
    .Y(_06476_));
 sky130_fd_sc_hd__nor2_1 _13740_ (.A(_05944_),
    .B(_06016_),
    .Y(_06477_));
 sky130_fd_sc_hd__or3_1 _13741_ (.A(_05946_),
    .B(_05899_),
    .C(_06007_),
    .X(_06478_));
 sky130_fd_sc_hd__xnor2_1 _13742_ (.A(_06475_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__a22o_1 _13743_ (.A1(_06475_),
    .A2(_06476_),
    .B1(_06477_),
    .B2(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__xor2_1 _13744_ (.A(_06474_),
    .B(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__a32o_1 _13745_ (.A1(_06471_),
    .A2(_06472_),
    .A3(_06481_),
    .B1(_06474_),
    .B2(_06480_),
    .X(_06482_));
 sky130_fd_sc_hd__nand2_1 _13746_ (.A(_06469_),
    .B(_06471_),
    .Y(_06483_));
 sky130_fd_sc_hd__o22a_1 _13747_ (.A1(_06065_),
    .A2(_06240_),
    .B1(_06161_),
    .B2(_05824_),
    .X(_06484_));
 sky130_fd_sc_hd__a21oi_1 _13748_ (.A1(_06383_),
    .A2(_06432_),
    .B1(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__xor2_1 _13749_ (.A(_06483_),
    .B(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__xor2_1 _13750_ (.A(_06468_),
    .B(_06482_),
    .X(_06487_));
 sky130_fd_sc_hd__nand2_1 _13751_ (.A(_06486_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__a21bo_1 _13752_ (.A1(_06468_),
    .A2(_06482_),
    .B1_N(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__and2b_1 _13753_ (.A_N(_06467_),
    .B(_06489_),
    .X(_06490_));
 sky130_fd_sc_hd__nand2_1 _13754_ (.A(_06483_),
    .B(_06485_),
    .Y(_06491_));
 sky130_fd_sc_hd__xor2_1 _13755_ (.A(_06467_),
    .B(_06489_),
    .X(_06492_));
 sky130_fd_sc_hd__nor2_1 _13756_ (.A(_06491_),
    .B(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__xor2_1 _13757_ (.A(_06438_),
    .B(_06455_),
    .X(_06494_));
 sky130_fd_sc_hd__o21ai_1 _13758_ (.A1(_06490_),
    .A2(_06493_),
    .B1(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__a211o_1 _13759_ (.A1(_06461_),
    .A2(_06458_),
    .B1(_06465_),
    .C1(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__nand3b_1 _13760_ (.A_N(_06426_),
    .B(_06462_),
    .C(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__a21bo_1 _13761_ (.A1(_06462_),
    .A2(_06496_),
    .B1_N(_06426_),
    .X(_06498_));
 sky130_fd_sc_hd__and3_1 _13762_ (.A(_06461_),
    .B(_06458_),
    .C(_06460_),
    .X(_06499_));
 sky130_fd_sc_hd__and2_1 _13763_ (.A(_06491_),
    .B(_06492_),
    .X(_06500_));
 sky130_fd_sc_hd__or4_1 _13764_ (.A(_06065_),
    .B(_05947_),
    .C(_05975_),
    .D(_05984_),
    .X(_06501_));
 sky130_fd_sc_hd__a2bb2o_1 _13765_ (.A1_N(_06065_),
    .A2_N(_06031_),
    .B1(_06002_),
    .B2(_05877_),
    .X(_06502_));
 sky130_fd_sc_hd__nand4_1 _13766_ (.A(_05855_),
    .B(_06153_),
    .C(_06501_),
    .D(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__and2_1 _13767_ (.A(_06501_),
    .B(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__or3_1 _13768_ (.A(_05825_),
    .B(_06240_),
    .C(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__or2_1 _13769_ (.A(_06486_),
    .B(_06487_),
    .X(_06506_));
 sky130_fd_sc_hd__and2_1 _13770_ (.A(_06488_),
    .B(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__nand2_1 _13771_ (.A(_06471_),
    .B(_06472_),
    .Y(_06508_));
 sky130_fd_sc_hd__xnor2_1 _13772_ (.A(_06508_),
    .B(_06481_),
    .Y(_06509_));
 sky130_fd_sc_hd__nor2_1 _13773_ (.A(_05823_),
    .B(_06045_),
    .Y(_06510_));
 sky130_fd_sc_hd__or3b_1 _13774_ (.A(_05944_),
    .B(_06009_),
    .C_N(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__o21bai_1 _13775_ (.A1(_06061_),
    .A2(_06009_),
    .B1_N(_06510_),
    .Y(_06512_));
 sky130_fd_sc_hd__a21bo_1 _13776_ (.A1(_06406_),
    .A2(_06511_),
    .B1_N(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__xor2_1 _13777_ (.A(_06477_),
    .B(_06479_),
    .X(_06514_));
 sky130_fd_sc_hd__and2b_1 _13778_ (.A_N(_06513_),
    .B(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__a22o_1 _13779_ (.A1(_05855_),
    .A2(_06153_),
    .B1(_06501_),
    .B2(_06502_),
    .X(_06516_));
 sky130_fd_sc_hd__xnor2_1 _13780_ (.A(_06514_),
    .B(_06513_),
    .Y(_06517_));
 sky130_fd_sc_hd__and3_1 _13781_ (.A(_06503_),
    .B(_06516_),
    .C(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__or2_1 _13782_ (.A(_06515_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__xnor2_1 _13783_ (.A(_06432_),
    .B(_06504_),
    .Y(_06520_));
 sky130_fd_sc_hd__xor2_1 _13784_ (.A(_06509_),
    .B(_06519_),
    .X(_06521_));
 sky130_fd_sc_hd__and2_1 _13785_ (.A(_06520_),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__a21o_1 _13786_ (.A1(_06509_),
    .A2(_06519_),
    .B1(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__nor2_1 _13787_ (.A(_06507_),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__nand2_1 _13788_ (.A(_06507_),
    .B(_06523_),
    .Y(_06525_));
 sky130_fd_sc_hd__nor2_1 _13789_ (.A(_06520_),
    .B(_06521_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand2_1 _13790_ (.A(_06382_),
    .B(_06002_),
    .Y(_06527_));
 sky130_fd_sc_hd__nor2_1 _13791_ (.A(_05824_),
    .B(_06031_),
    .Y(_06528_));
 sky130_fd_sc_hd__xnor2_1 _13792_ (.A(_06527_),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__nand2_1 _13793_ (.A(_05855_),
    .B(_06061_),
    .Y(_06530_));
 sky130_fd_sc_hd__nand2_1 _13794_ (.A(_06511_),
    .B(_06512_),
    .Y(_06531_));
 sky130_fd_sc_hd__o21ba_1 _13795_ (.A1(_06057_),
    .A2(_06530_),
    .B1_N(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__a41o_1 _13796_ (.A1(_05855_),
    .A2(_05877_),
    .A3(_06061_),
    .A4(_06078_),
    .B1(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__nand2_1 _13797_ (.A(_06529_),
    .B(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__nor2_1 _13798_ (.A(_05877_),
    .B(_05888_),
    .Y(_06535_));
 sky130_fd_sc_hd__nor2_1 _13799_ (.A(_06057_),
    .B(_06061_),
    .Y(_06536_));
 sky130_fd_sc_hd__nor2_1 _13800_ (.A(_06529_),
    .B(_06533_),
    .Y(_06537_));
 sky130_fd_sc_hd__or4_1 _13801_ (.A(_05824_),
    .B(_06535_),
    .C(_06536_),
    .D(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__nand3b_1 _13802_ (.A_N(_06406_),
    .B(_06531_),
    .C(_06530_),
    .Y(_06539_));
 sky130_fd_sc_hd__a21oi_1 _13803_ (.A1(_06503_),
    .A2(_06516_),
    .B1(_06517_),
    .Y(_06540_));
 sky130_fd_sc_hd__a311o_1 _13804_ (.A1(_06534_),
    .A2(_06538_),
    .A3(_06539_),
    .B1(_06540_),
    .C1(_06518_),
    .X(_06541_));
 sky130_fd_sc_hd__o31a_1 _13805_ (.A1(_05825_),
    .A2(_06031_),
    .A3(_06527_),
    .B1(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__or4_1 _13806_ (.A(_06522_),
    .B(_06524_),
    .C(_06526_),
    .D(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__o211a_1 _13807_ (.A1(_06505_),
    .A2(_06524_),
    .B1(_06525_),
    .C1(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__or3_1 _13808_ (.A(_06490_),
    .B(_06493_),
    .C(_06494_),
    .X(_06545_));
 sky130_fd_sc_hd__or4b_1 _13809_ (.A(_06500_),
    .B(_06493_),
    .C(_06544_),
    .D_N(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__or3_1 _13810_ (.A(_06499_),
    .B(_06465_),
    .C(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__a21oi_1 _13811_ (.A1(_06497_),
    .A2(_06498_),
    .B1(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__nor2_1 _13812_ (.A(_06426_),
    .B(_06496_),
    .Y(_06549_));
 sky130_fd_sc_hd__o21bai_1 _13813_ (.A1(_06426_),
    .A2(_06462_),
    .B1_N(_06422_),
    .Y(_06550_));
 sky130_fd_sc_hd__xor2_1 _13814_ (.A(_06423_),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__o21ai_1 _13815_ (.A1(_06548_),
    .A2(_06549_),
    .B1(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__o21ba_1 _13816_ (.A1(_06336_),
    .A2(_06375_),
    .B1_N(_06424_),
    .X(_06553_));
 sky130_fd_sc_hd__xor2_1 _13817_ (.A(_06376_),
    .B(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__a21bo_1 _13818_ (.A1(_06464_),
    .A2(_06552_),
    .B1_N(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__nor2_1 _13819_ (.A(_06333_),
    .B(_06377_),
    .Y(_06556_));
 sky130_fd_sc_hd__xnor2_2 _13820_ (.A(_06279_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__a21bo_1 _13821_ (.A1(_06425_),
    .A2(_06555_),
    .B1_N(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__xnor2_1 _13822_ (.A(_06278_),
    .B(_06334_),
    .Y(_06559_));
 sky130_fd_sc_hd__a21o_2 _13823_ (.A1(_06378_),
    .A2(_06558_),
    .B1(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(_06193_),
    .B(_06231_),
    .Y(_06561_));
 sky130_fd_sc_hd__xor2_2 _13825_ (.A(_06561_),
    .B(_06276_),
    .X(_06562_));
 sky130_fd_sc_hd__a21oi_4 _13826_ (.A1(_06335_),
    .A2(_06560_),
    .B1(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__and2_1 _13827_ (.A(_06232_),
    .B(_06275_),
    .X(_06564_));
 sky130_fd_sc_hd__or2b_1 _13828_ (.A(_06268_),
    .B_N(_06235_),
    .X(_06565_));
 sky130_fd_sc_hd__or2b_1 _13829_ (.A(_06271_),
    .B_N(_06269_),
    .X(_06566_));
 sky130_fd_sc_hd__nand2_1 _13830_ (.A(_06565_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__a21bo_1 _13831_ (.A1(_06253_),
    .A2(_06267_),
    .B1_N(_06251_),
    .X(_06568_));
 sky130_fd_sc_hd__or3_1 _13832_ (.A(_05974_),
    .B(_06161_),
    .C(_05940_),
    .X(_06569_));
 sky130_fd_sc_hd__o21ai_1 _13833_ (.A1(_05974_),
    .A2(_06245_),
    .B1(_06161_),
    .Y(_06570_));
 sky130_fd_sc_hd__nand2_1 _13834_ (.A(_06569_),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__a21o_1 _13835_ (.A1(_06242_),
    .A2(_06244_),
    .B1(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__nand3_1 _13836_ (.A(_06242_),
    .B(_06244_),
    .C(_06571_),
    .Y(_06573_));
 sky130_fd_sc_hd__and2_1 _13837_ (.A(_06572_),
    .B(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__and2b_1 _13838_ (.A_N(_06258_),
    .B(_06261_),
    .X(_06575_));
 sky130_fd_sc_hd__or4_1 _13839_ (.A(_06015_),
    .B(_05991_),
    .C(_05978_),
    .D(_06055_),
    .X(_06576_));
 sky130_fd_sc_hd__a32o_1 _13840_ (.A1(_05752_),
    .A2(_05921_),
    .A3(_06053_),
    .B1(_05974_),
    .B2(_05989_),
    .X(_06577_));
 sky130_fd_sc_hd__and2_1 _13841_ (.A(_06576_),
    .B(_06577_),
    .X(_06578_));
 sky130_fd_sc_hd__o21ai_1 _13842_ (.A1(_06259_),
    .A2(_06575_),
    .B1(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__or3_1 _13843_ (.A(_06259_),
    .B(_06575_),
    .C(_06578_),
    .X(_06580_));
 sky130_fd_sc_hd__and2_1 _13844_ (.A(_06579_),
    .B(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__xnor2_1 _13845_ (.A(_06248_),
    .B(_06581_),
    .Y(_06582_));
 sky130_fd_sc_hd__nor2_1 _13846_ (.A(_06263_),
    .B(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__and2_1 _13847_ (.A(_06263_),
    .B(_06582_),
    .X(_06584_));
 sky130_fd_sc_hd__nor2_1 _13848_ (.A(_06583_),
    .B(_06584_),
    .Y(_06585_));
 sky130_fd_sc_hd__nand2_1 _13849_ (.A(_06574_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__or2_1 _13850_ (.A(_06574_),
    .B(_06585_),
    .X(_06587_));
 sky130_fd_sc_hd__nand2_1 _13851_ (.A(_06586_),
    .B(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__xnor2_1 _13852_ (.A(_06568_),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__nor2_1 _13853_ (.A(_06219_),
    .B(_06266_),
    .Y(_06590_));
 sky130_fd_sc_hd__a21oi_1 _13854_ (.A1(_06255_),
    .A2(_06265_),
    .B1(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__xor2_1 _13855_ (.A(_06589_),
    .B(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__xnor2_1 _13856_ (.A(_06567_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__xor2_1 _13857_ (.A(_06273_),
    .B(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__nand2_2 _13858_ (.A(_06564_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__or2_1 _13859_ (.A(_06564_),
    .B(_06594_),
    .X(_06596_));
 sky130_fd_sc_hd__nand2_1 _13860_ (.A(_06595_),
    .B(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__o21bai_4 _13861_ (.A1(_06277_),
    .A2(_06563_),
    .B1_N(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__or3b_1 _13862_ (.A(_06277_),
    .B(_06563_),
    .C_N(_06597_),
    .X(_06599_));
 sky130_fd_sc_hd__and3_1 _13863_ (.A(_06335_),
    .B(_06560_),
    .C(_06562_),
    .X(_06600_));
 sky130_fd_sc_hd__nand3_1 _13864_ (.A(_06559_),
    .B(_06378_),
    .C(_06558_),
    .Y(_06601_));
 sky130_fd_sc_hd__nand2_2 _13865_ (.A(_06425_),
    .B(_06555_),
    .Y(_06602_));
 sky130_fd_sc_hd__xor2_4 _13866_ (.A(_06602_),
    .B(_06557_),
    .X(_06603_));
 sky130_fd_sc_hd__nand2_1 _13867_ (.A(_06464_),
    .B(_06552_),
    .Y(_06604_));
 sky130_fd_sc_hd__xnor2_2 _13868_ (.A(_06604_),
    .B(_06554_),
    .Y(_06605_));
 sky130_fd_sc_hd__or3_1 _13869_ (.A(_06548_),
    .B(_06549_),
    .C(_06551_),
    .X(_06606_));
 sky130_fd_sc_hd__and2_2 _13870_ (.A(_06552_),
    .B(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__and3_1 _13871_ (.A(_06547_),
    .B(_06497_),
    .C(_06498_),
    .X(_06608_));
 sky130_fd_sc_hd__or2_1 _13872_ (.A(_06548_),
    .B(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__clkbuf_4 _13873_ (.A(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__and2b_1 _13874_ (.A_N(_06607_),
    .B(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__nor2_4 _13875_ (.A(_06605_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__a211oi_2 _13876_ (.A1(_06560_),
    .A2(_06601_),
    .B1(_06603_),
    .C1(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__o21ai_2 _13877_ (.A1(_06563_),
    .A2(_06600_),
    .B1(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__a21oi_4 _13878_ (.A1(_06598_),
    .A2(_06599_),
    .B1(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_1 _13879_ (.A(_06273_),
    .B(_06593_),
    .Y(_06616_));
 sky130_fd_sc_hd__and2b_1 _13880_ (.A_N(_06592_),
    .B(_06567_),
    .X(_06617_));
 sky130_fd_sc_hd__and2b_1 _13881_ (.A_N(_06591_),
    .B(_06589_),
    .X(_06618_));
 sky130_fd_sc_hd__a31o_1 _13882_ (.A1(_06568_),
    .A2(_06586_),
    .A3(_06587_),
    .B1(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__or3_1 _13883_ (.A(_06239_),
    .B(_06245_),
    .C(_06202_),
    .X(_06620_));
 sky130_fd_sc_hd__nor2_1 _13884_ (.A(_06201_),
    .B(_06052_),
    .Y(_06621_));
 sky130_fd_sc_hd__or2_1 _13885_ (.A(_05978_),
    .B(_06067_),
    .X(_06622_));
 sky130_fd_sc_hd__nand2_1 _13886_ (.A(_05974_),
    .B(_05983_),
    .Y(_06623_));
 sky130_fd_sc_hd__and3_1 _13887_ (.A(_06201_),
    .B(_06052_),
    .C(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__xnor2_1 _13888_ (.A(_06622_),
    .B(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__o21a_1 _13889_ (.A1(_06621_),
    .A2(_06625_),
    .B1(_06576_),
    .X(_06626_));
 sky130_fd_sc_hd__inv_2 _13890_ (.A(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__xnor2_1 _13891_ (.A(_06572_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__or2_1 _13892_ (.A(_06579_),
    .B(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__nand2_1 _13893_ (.A(_06579_),
    .B(_06628_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand2_1 _13894_ (.A(_06629_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__or2_1 _13895_ (.A(_06620_),
    .B(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__nand2_1 _13896_ (.A(_06620_),
    .B(_06631_),
    .Y(_06633_));
 sky130_fd_sc_hd__and2_1 _13897_ (.A(_06632_),
    .B(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__xnor2_2 _13898_ (.A(_06586_),
    .B(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__a21o_1 _13899_ (.A1(_06248_),
    .A2(_06581_),
    .B1(_06583_),
    .X(_06636_));
 sky130_fd_sc_hd__xnor2_2 _13900_ (.A(_06635_),
    .B(_06636_),
    .Y(_06637_));
 sky130_fd_sc_hd__xnor2_2 _13901_ (.A(_06619_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__xor2_2 _13902_ (.A(_06617_),
    .B(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__xnor2_2 _13903_ (.A(_06616_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__nand3_4 _13904_ (.A(_06595_),
    .B(_06598_),
    .C(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__a21o_2 _13905_ (.A1(_06595_),
    .A2(_06598_),
    .B1(_06640_),
    .X(_06642_));
 sky130_fd_sc_hd__inv_2 _13906_ (.A(_06640_),
    .Y(_06643_));
 sky130_fd_sc_hd__and2b_1 _13907_ (.A_N(_06637_),
    .B(_06619_),
    .X(_06644_));
 sky130_fd_sc_hd__a32o_1 _13908_ (.A1(_06574_),
    .A2(_06585_),
    .A3(_06634_),
    .B1(_06635_),
    .B2(_06636_),
    .X(_06645_));
 sky130_fd_sc_hd__a21oi_1 _13909_ (.A1(_05752_),
    .A2(_06201_),
    .B1(_06621_),
    .Y(_06646_));
 sky130_fd_sc_hd__a41o_1 _13910_ (.A1(_05752_),
    .A2(_05989_),
    .A3(_06053_),
    .A4(_06624_),
    .B1(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__xnor2_1 _13911_ (.A(_06569_),
    .B(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__nand2_1 _13912_ (.A(_06576_),
    .B(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__xnor2_1 _13913_ (.A(_06632_),
    .B(_06649_),
    .Y(_06650_));
 sky130_fd_sc_hd__o211a_1 _13914_ (.A1(_06572_),
    .A2(_06627_),
    .B1(_06629_),
    .C1(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__xnor2_1 _13915_ (.A(_06645_),
    .B(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__xnor2_1 _13916_ (.A(_06644_),
    .B(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(_06616_),
    .B(_06595_),
    .Y(_06654_));
 sky130_fd_sc_hd__and2_1 _13918_ (.A(_06617_),
    .B(_06638_),
    .X(_06655_));
 sky130_fd_sc_hd__a21oi_1 _13919_ (.A1(_06639_),
    .A2(_06654_),
    .B1(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__o211a_1 _13920_ (.A1(_06598_),
    .A2(_06643_),
    .B1(_06653_),
    .C1(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__a31o_4 _13921_ (.A1(_06615_),
    .A2(_06641_),
    .A3(_06642_),
    .B1(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__nor2_2 _13922_ (.A(_05825_),
    .B(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__o211a_1 _13923_ (.A1(_06603_),
    .A2(_06612_),
    .B1(_06560_),
    .C1(_06601_),
    .X(_06660_));
 sky130_fd_sc_hd__or2_1 _13924_ (.A(_06613_),
    .B(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__clkbuf_2 _13925_ (.A(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_4 _13926_ (.A(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__nor2_2 _13927_ (.A(_06031_),
    .B(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand2_1 _13928_ (.A(_06659_),
    .B(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__clkbuf_4 _13929_ (.A(_05982_),
    .X(_06666_));
 sky130_fd_sc_hd__xnor2_4 _13930_ (.A(_06603_),
    .B(_06612_),
    .Y(_06667_));
 sky130_fd_sc_hd__clkbuf_4 _13931_ (.A(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__xnor2_1 _13932_ (.A(_06659_),
    .B(_06664_),
    .Y(_06669_));
 sky130_fd_sc_hd__or3_1 _13933_ (.A(_06666_),
    .B(_06668_),
    .C(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__xor2_4 _13934_ (.A(_06607_),
    .B(_06610_),
    .X(_06671_));
 sky130_fd_sc_hd__clkbuf_4 _13935_ (.A(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__nor2_1 _13936_ (.A(_06245_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nor2_2 _13937_ (.A(_06161_),
    .B(_06667_),
    .Y(_06674_));
 sky130_fd_sc_hd__clkbuf_4 _13938_ (.A(_06240_),
    .X(_06675_));
 sky130_fd_sc_hd__and2_1 _13939_ (.A(_06605_),
    .B(_06611_),
    .X(_06676_));
 sky130_fd_sc_hd__nor2_4 _13940_ (.A(_06612_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__clkbuf_4 _13941_ (.A(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__nor2_1 _13942_ (.A(_06675_),
    .B(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__clkbuf_4 _13943_ (.A(_06161_),
    .X(_06680_));
 sky130_fd_sc_hd__nor2_1 _13944_ (.A(_06680_),
    .B(_06677_),
    .Y(_06681_));
 sky130_fd_sc_hd__o21ba_1 _13945_ (.A1(_06675_),
    .A2(_06668_),
    .B1_N(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a21oi_1 _13946_ (.A1(_06674_),
    .A2(_06679_),
    .B1(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__xnor2_1 _13947_ (.A(_06673_),
    .B(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__a21o_1 _13948_ (.A1(_06665_),
    .A2(_06670_),
    .B1(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__nand3_1 _13949_ (.A(_06665_),
    .B(_06670_),
    .C(_06684_),
    .Y(_06686_));
 sky130_fd_sc_hd__nand2_1 _13950_ (.A(_06685_),
    .B(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__nor2_1 _13951_ (.A(_06675_),
    .B(_06672_),
    .Y(_06688_));
 sky130_fd_sc_hd__clkbuf_4 _13952_ (.A(_06245_),
    .X(_06689_));
 sky130_fd_sc_hd__clkbuf_4 _13953_ (.A(_06610_),
    .X(_06690_));
 sky130_fd_sc_hd__or2_1 _13954_ (.A(_06689_),
    .B(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__nor2_1 _13955_ (.A(_06680_),
    .B(_06672_),
    .Y(_06692_));
 sky130_fd_sc_hd__nor2_1 _13956_ (.A(_06679_),
    .B(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__o2bb2a_1 _13957_ (.A1_N(_06681_),
    .A2_N(_06688_),
    .B1(_06691_),
    .B2(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__or2_1 _13958_ (.A(_06687_),
    .B(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__clkbuf_4 _13959_ (.A(_06080_),
    .X(_06696_));
 sky130_fd_sc_hd__nor2_1 _13960_ (.A(_06696_),
    .B(_06671_),
    .Y(_06697_));
 sky130_fd_sc_hd__clkbuf_4 _13961_ (.A(_06134_),
    .X(_06698_));
 sky130_fd_sc_hd__nor2_2 _13962_ (.A(_06698_),
    .B(_06690_),
    .Y(_06699_));
 sky130_fd_sc_hd__nand2_2 _13963_ (.A(_06697_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__o22ai_1 _13964_ (.A1(_06696_),
    .A2(_06690_),
    .B1(_06672_),
    .B2(_06698_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand2_1 _13965_ (.A(_06700_),
    .B(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__a21oi_2 _13966_ (.A1(_06685_),
    .A2(_06695_),
    .B1(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__clkbuf_4 _13967_ (.A(_06031_),
    .X(_06704_));
 sky130_fd_sc_hd__nor2_2 _13968_ (.A(_06704_),
    .B(_06658_),
    .Y(_06705_));
 sky130_fd_sc_hd__or3_1 _13969_ (.A(_06613_),
    .B(_06563_),
    .C(_06600_),
    .X(_06706_));
 sky130_fd_sc_hd__nand2_2 _13970_ (.A(_06614_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__clkbuf_4 _13971_ (.A(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__nor2_1 _13972_ (.A(_05825_),
    .B(_06708_),
    .Y(_06709_));
 sky130_fd_sc_hd__nand2_1 _13973_ (.A(_06705_),
    .B(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__nor2_1 _13974_ (.A(_06031_),
    .B(_06707_),
    .Y(_06711_));
 sky130_fd_sc_hd__xnor2_1 _13975_ (.A(_06659_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__or3_1 _13976_ (.A(_05982_),
    .B(_06663_),
    .C(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__or2_1 _13977_ (.A(_06240_),
    .B(_06662_),
    .X(_06714_));
 sky130_fd_sc_hd__xnor2_1 _13978_ (.A(_06714_),
    .B(_06674_),
    .Y(_06715_));
 sky130_fd_sc_hd__or3b_1 _13979_ (.A(_06245_),
    .B(_06678_),
    .C_N(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__o21bai_1 _13980_ (.A1(_06245_),
    .A2(_06678_),
    .B1_N(_06715_),
    .Y(_06717_));
 sky130_fd_sc_hd__nand2_1 _13981_ (.A(_06716_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__a21o_1 _13982_ (.A1(_06710_),
    .A2(_06713_),
    .B1(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__a22oi_2 _13983_ (.A1(_06674_),
    .A2(_06679_),
    .B1(_06673_),
    .B2(_06683_),
    .Y(_06720_));
 sky130_fd_sc_hd__nand3_1 _13984_ (.A(_06710_),
    .B(_06713_),
    .C(_06718_),
    .Y(_06721_));
 sky130_fd_sc_hd__and2_1 _13985_ (.A(_06719_),
    .B(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__or2b_1 _13986_ (.A(_06720_),
    .B_N(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__clkbuf_4 _13987_ (.A(_06067_),
    .X(_06724_));
 sky130_fd_sc_hd__nor2_1 _13988_ (.A(_06696_),
    .B(_06677_),
    .Y(_06725_));
 sky130_fd_sc_hd__inv_2 _13989_ (.A(_06725_),
    .Y(_06726_));
 sky130_fd_sc_hd__o21bai_1 _13990_ (.A1(_06134_),
    .A2(_06677_),
    .B1_N(_06697_),
    .Y(_06727_));
 sky130_fd_sc_hd__o31a_1 _13991_ (.A1(_06698_),
    .A2(_06726_),
    .A3(_06671_),
    .B1(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__or3b_1 _13992_ (.A(_06724_),
    .B(_06610_),
    .C_N(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__o21bai_1 _13993_ (.A1(_06724_),
    .A2(_06690_),
    .B1_N(_06728_),
    .Y(_06730_));
 sky130_fd_sc_hd__nand2_1 _13994_ (.A(_06729_),
    .B(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__nor2_1 _13995_ (.A(_06731_),
    .B(_06700_),
    .Y(_06732_));
 sky130_fd_sc_hd__and2_1 _13996_ (.A(_06731_),
    .B(_06700_),
    .X(_06733_));
 sky130_fd_sc_hd__or2_1 _13997_ (.A(_06732_),
    .B(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__a21oi_2 _13998_ (.A1(_06719_),
    .A2(_06723_),
    .B1(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__and3_1 _13999_ (.A(_06719_),
    .B(_06723_),
    .C(_06734_),
    .X(_06736_));
 sky130_fd_sc_hd__nor2_1 _14000_ (.A(_06735_),
    .B(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__and3_1 _14001_ (.A(_06614_),
    .B(_06598_),
    .C(_06599_),
    .X(_06738_));
 sky130_fd_sc_hd__or2_1 _14002_ (.A(_06615_),
    .B(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__clkbuf_4 _14003_ (.A(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__nor2_1 _14004_ (.A(_06704_),
    .B(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__xnor2_1 _14005_ (.A(_06659_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _14006_ (.A(_06659_),
    .B(_06741_),
    .Y(_06743_));
 sky130_fd_sc_hd__o31ai_2 _14007_ (.A1(_06666_),
    .A2(_06708_),
    .A3(_06742_),
    .B1(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__nor2_1 _14008_ (.A(_06245_),
    .B(_06668_),
    .Y(_06745_));
 sky130_fd_sc_hd__nor2_1 _14009_ (.A(_06240_),
    .B(_06707_),
    .Y(_06746_));
 sky130_fd_sc_hd__nor2_1 _14010_ (.A(_06680_),
    .B(_06662_),
    .Y(_06747_));
 sky130_fd_sc_hd__nand2_1 _14011_ (.A(_06746_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__or2_1 _14012_ (.A(_06746_),
    .B(_06747_),
    .X(_06749_));
 sky130_fd_sc_hd__nand2_1 _14013_ (.A(_06748_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__xnor2_2 _14014_ (.A(_06745_),
    .B(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__xnor2_1 _14015_ (.A(_06744_),
    .B(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__o31ai_1 _14016_ (.A1(_06680_),
    .A2(_06668_),
    .A3(_06714_),
    .B1(_06716_),
    .Y(_06753_));
 sky130_fd_sc_hd__inv_2 _14017_ (.A(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__nor2_1 _14018_ (.A(_06752_),
    .B(_06754_),
    .Y(_06755_));
 sky130_fd_sc_hd__and2_1 _14019_ (.A(_06752_),
    .B(_06754_),
    .X(_06756_));
 sky130_fd_sc_hd__nor2_1 _14020_ (.A(_06755_),
    .B(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand3_4 _14021_ (.A(_06615_),
    .B(_06641_),
    .C(_06642_),
    .Y(_06758_));
 sky130_fd_sc_hd__a21o_2 _14022_ (.A1(_06641_),
    .A2(_06642_),
    .B1(_06615_),
    .X(_06759_));
 sky130_fd_sc_hd__nand2_4 _14023_ (.A(_06758_),
    .B(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_2 _14024_ (.A(_05752_),
    .B(_06658_),
    .Y(_06761_));
 sky130_fd_sc_hd__o22ai_2 _14025_ (.A1(_06704_),
    .A2(_06760_),
    .B1(_06761_),
    .B2(_05825_),
    .Y(_06762_));
 sky130_fd_sc_hd__nand3_2 _14026_ (.A(_05855_),
    .B(_06758_),
    .C(_06759_),
    .Y(_06763_));
 sky130_fd_sc_hd__or3_1 _14027_ (.A(_06704_),
    .B(_06761_),
    .C(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__nor2_1 _14028_ (.A(_05982_),
    .B(_06740_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand3_1 _14029_ (.A(_06762_),
    .B(_06764_),
    .C(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__a21o_1 _14030_ (.A1(_06762_),
    .A2(_06764_),
    .B1(_06765_),
    .X(_06767_));
 sky130_fd_sc_hd__nand2_1 _14031_ (.A(_06766_),
    .B(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__clkbuf_4 _14032_ (.A(_06016_),
    .X(_06769_));
 sky130_fd_sc_hd__a311oi_4 _14033_ (.A1(_06615_),
    .A2(_06641_),
    .A3(_06642_),
    .B1(_06657_),
    .C1(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__and2_1 _14034_ (.A(_06002_),
    .B(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a21o_1 _14035_ (.A1(_05984_),
    .A2(_06769_),
    .B1(_06658_),
    .X(_06772_));
 sky130_fd_sc_hd__nor2_1 _14036_ (.A(_06009_),
    .B(_06658_),
    .Y(_06773_));
 sky130_fd_sc_hd__or3b_1 _14037_ (.A(_06771_),
    .B(_06772_),
    .C_N(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__o21bai_1 _14038_ (.A1(_06771_),
    .A2(_06772_),
    .B1_N(_06773_),
    .Y(_06775_));
 sky130_fd_sc_hd__buf_2 _14039_ (.A(_05984_),
    .X(_06776_));
 sky130_fd_sc_hd__nor2_1 _14040_ (.A(_06776_),
    .B(_06658_),
    .Y(_06777_));
 sky130_fd_sc_hd__and3_1 _14041_ (.A(_06012_),
    .B(_06758_),
    .C(_06759_),
    .X(_06778_));
 sky130_fd_sc_hd__a31o_1 _14042_ (.A1(_06002_),
    .A2(_06758_),
    .A3(_06759_),
    .B1(_06770_),
    .X(_06779_));
 sky130_fd_sc_hd__a22o_1 _14043_ (.A1(_06777_),
    .A2(_06778_),
    .B1(_06779_),
    .B2(_06773_),
    .X(_06780_));
 sky130_fd_sc_hd__and3_1 _14044_ (.A(_06774_),
    .B(_06775_),
    .C(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__a21o_1 _14045_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06780_),
    .X(_06782_));
 sky130_fd_sc_hd__or2b_1 _14046_ (.A(_06781_),
    .B_N(_06782_),
    .X(_06783_));
 sky130_fd_sc_hd__xnor2_1 _14047_ (.A(_06768_),
    .B(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__nor2_1 _14048_ (.A(_06666_),
    .B(_06708_),
    .Y(_06785_));
 sky130_fd_sc_hd__xnor2_1 _14049_ (.A(_06742_),
    .B(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__inv_2 _14050_ (.A(_06773_),
    .Y(_06787_));
 sky130_fd_sc_hd__a21bo_1 _14051_ (.A1(_06777_),
    .A2(_06778_),
    .B1_N(_06779_),
    .X(_06788_));
 sky130_fd_sc_hd__xnor2_1 _14052_ (.A(_06787_),
    .B(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__nor2_1 _14053_ (.A(_06776_),
    .B(_06739_),
    .Y(_06790_));
 sky130_fd_sc_hd__xnor2_1 _14054_ (.A(_06778_),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__nand2_1 _14055_ (.A(_06778_),
    .B(_06790_),
    .Y(_06792_));
 sky130_fd_sc_hd__o21ai_1 _14056_ (.A1(_06787_),
    .A2(_06791_),
    .B1(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__xnor2_1 _14057_ (.A(_06789_),
    .B(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__or2b_1 _14058_ (.A(_06789_),
    .B_N(_06793_),
    .X(_06795_));
 sky130_fd_sc_hd__a21bo_1 _14059_ (.A1(_06786_),
    .A2(_06794_),
    .B1_N(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__xnor2_1 _14060_ (.A(_06784_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__xnor2_1 _14061_ (.A(_06757_),
    .B(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__xnor2_1 _14062_ (.A(_06722_),
    .B(_06720_),
    .Y(_06799_));
 sky130_fd_sc_hd__xor2_1 _14063_ (.A(_06786_),
    .B(_06794_),
    .X(_06800_));
 sky130_fd_sc_hd__o21ai_1 _14064_ (.A1(_06666_),
    .A2(_06663_),
    .B1(_06712_),
    .Y(_06801_));
 sky130_fd_sc_hd__and2_1 _14065_ (.A(_06713_),
    .B(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__xnor2_1 _14066_ (.A(_06787_),
    .B(_06791_),
    .Y(_06803_));
 sky130_fd_sc_hd__or2_1 _14067_ (.A(_06769_),
    .B(_06707_),
    .X(_06804_));
 sky130_fd_sc_hd__buf_2 _14068_ (.A(_06009_),
    .X(_06805_));
 sky130_fd_sc_hd__and3b_1 _14069_ (.A_N(_06805_),
    .B(_06758_),
    .C(_06759_),
    .X(_06806_));
 sky130_fd_sc_hd__o32ai_1 _14070_ (.A1(_06769_),
    .A2(_06615_),
    .A3(_06738_),
    .B1(_06707_),
    .B2(_06776_),
    .Y(_06807_));
 sky130_fd_sc_hd__o31a_1 _14071_ (.A1(_06776_),
    .A2(_06739_),
    .A3(_06804_),
    .B1(_06807_),
    .X(_06808_));
 sky130_fd_sc_hd__nand2_1 _14072_ (.A(_06806_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__o31a_1 _14073_ (.A1(_06776_),
    .A2(_06740_),
    .A3(_06804_),
    .B1(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__xor2_1 _14074_ (.A(_06803_),
    .B(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__nor2_1 _14075_ (.A(_06803_),
    .B(_06810_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21oi_1 _14076_ (.A1(_06802_),
    .A2(_06811_),
    .B1(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__xnor2_1 _14077_ (.A(_06800_),
    .B(_06813_),
    .Y(_06814_));
 sky130_fd_sc_hd__or2b_1 _14078_ (.A(_06813_),
    .B_N(_06800_),
    .X(_06815_));
 sky130_fd_sc_hd__a21bo_1 _14079_ (.A1(_06799_),
    .A2(_06814_),
    .B1_N(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__xnor2_2 _14080_ (.A(_06798_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__xnor2_2 _14081_ (.A(_06737_),
    .B(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__and3_1 _14082_ (.A(_06685_),
    .B(_06695_),
    .C(_06702_),
    .X(_06819_));
 sky130_fd_sc_hd__nor2_1 _14083_ (.A(_06703_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__xnor2_1 _14084_ (.A(_06799_),
    .B(_06814_),
    .Y(_06821_));
 sky130_fd_sc_hd__xor2_1 _14085_ (.A(_06687_),
    .B(_06694_),
    .X(_06822_));
 sky130_fd_sc_hd__xnor2_1 _14086_ (.A(_06802_),
    .B(_06811_),
    .Y(_06823_));
 sky130_fd_sc_hd__nor2_1 _14087_ (.A(_06666_),
    .B(_06668_),
    .Y(_06824_));
 sky130_fd_sc_hd__xnor2_1 _14088_ (.A(_06669_),
    .B(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__xnor2_1 _14089_ (.A(_06806_),
    .B(_06808_),
    .Y(_06826_));
 sky130_fd_sc_hd__nor2_1 _14090_ (.A(_06805_),
    .B(_06740_),
    .Y(_06827_));
 sky130_fd_sc_hd__nor2_1 _14091_ (.A(_06776_),
    .B(_06662_),
    .Y(_06828_));
 sky130_fd_sc_hd__xnor2_1 _14092_ (.A(_06804_),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__and2b_1 _14093_ (.A_N(_06804_),
    .B(_06828_),
    .X(_06830_));
 sky130_fd_sc_hd__a21oi_1 _14094_ (.A1(_06827_),
    .A2(_06829_),
    .B1(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__xor2_1 _14095_ (.A(_06826_),
    .B(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__nor2_1 _14096_ (.A(_06826_),
    .B(_06831_),
    .Y(_06833_));
 sky130_fd_sc_hd__a21o_1 _14097_ (.A1(_06825_),
    .A2(_06832_),
    .B1(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__xnor2_1 _14098_ (.A(_06823_),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__or2b_1 _14099_ (.A(_06823_),
    .B_N(_06834_),
    .X(_06836_));
 sky130_fd_sc_hd__a21boi_1 _14100_ (.A1(_06822_),
    .A2(_06835_),
    .B1_N(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__xor2_1 _14101_ (.A(_06821_),
    .B(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__nor2_1 _14102_ (.A(_06821_),
    .B(_06837_),
    .Y(_06839_));
 sky130_fd_sc_hd__a21oi_2 _14103_ (.A1(_06820_),
    .A2(_06838_),
    .B1(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__xor2_2 _14104_ (.A(_06818_),
    .B(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__xnor2_2 _14105_ (.A(_06703_),
    .B(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__nor2_1 _14106_ (.A(_06704_),
    .B(_06760_),
    .Y(_06843_));
 sky130_fd_sc_hd__nor2_1 _14107_ (.A(_05825_),
    .B(_06668_),
    .Y(_06844_));
 sky130_fd_sc_hd__nor2_1 _14108_ (.A(_06704_),
    .B(_06668_),
    .Y(_06845_));
 sky130_fd_sc_hd__xnor2_2 _14109_ (.A(_06763_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__nor2_1 _14110_ (.A(_06666_),
    .B(_06678_),
    .Y(_06847_));
 sky130_fd_sc_hd__a22o_1 _14111_ (.A1(_06843_),
    .A2(_06844_),
    .B1(_06846_),
    .B2(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__a21oi_1 _14112_ (.A1(_06681_),
    .A2(_06688_),
    .B1(_06693_),
    .Y(_06849_));
 sky130_fd_sc_hd__xnor2_1 _14113_ (.A(_06691_),
    .B(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__xnor2_1 _14114_ (.A(_06848_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__nor2_1 _14115_ (.A(_06675_),
    .B(_06690_),
    .Y(_06852_));
 sky130_fd_sc_hd__and2_1 _14116_ (.A(_06692_),
    .B(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__and2b_1 _14117_ (.A_N(_06851_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__a21oi_1 _14118_ (.A1(_06848_),
    .A2(_06850_),
    .B1(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__and2b_1 _14119_ (.A_N(_06855_),
    .B(_06699_),
    .X(_06856_));
 sky130_fd_sc_hd__xnor2_1 _14120_ (.A(_06820_),
    .B(_06838_),
    .Y(_06857_));
 sky130_fd_sc_hd__xnor2_1 _14121_ (.A(_06699_),
    .B(_06855_),
    .Y(_06858_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_06822_),
    .B(_06835_),
    .Y(_06859_));
 sky130_fd_sc_hd__xnor2_1 _14123_ (.A(_06851_),
    .B(_06853_),
    .Y(_06860_));
 sky130_fd_sc_hd__xnor2_1 _14124_ (.A(_06825_),
    .B(_06832_),
    .Y(_06861_));
 sky130_fd_sc_hd__xor2_2 _14125_ (.A(_06846_),
    .B(_06847_),
    .X(_06862_));
 sky130_fd_sc_hd__xnor2_1 _14126_ (.A(_06827_),
    .B(_06829_),
    .Y(_06863_));
 sky130_fd_sc_hd__nor2_1 _14127_ (.A(_06769_),
    .B(_06667_),
    .Y(_06864_));
 sky130_fd_sc_hd__or2_1 _14128_ (.A(_06805_),
    .B(_06707_),
    .X(_06865_));
 sky130_fd_sc_hd__o22a_1 _14129_ (.A1(_06769_),
    .A2(_06662_),
    .B1(_06667_),
    .B2(_06776_),
    .X(_06866_));
 sky130_fd_sc_hd__a21o_1 _14130_ (.A1(_06828_),
    .A2(_06864_),
    .B1(_06866_),
    .X(_06867_));
 sky130_fd_sc_hd__o2bb2ai_1 _14131_ (.A1_N(_06828_),
    .A2_N(_06864_),
    .B1(_06865_),
    .B2(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__xnor2_1 _14132_ (.A(_06863_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__or2b_1 _14133_ (.A(_06863_),
    .B_N(_06868_),
    .X(_06870_));
 sky130_fd_sc_hd__a21boi_1 _14134_ (.A1(_06862_),
    .A2(_06869_),
    .B1_N(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__nor2_1 _14135_ (.A(_06861_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__nand2_1 _14136_ (.A(_06861_),
    .B(_06871_),
    .Y(_06873_));
 sky130_fd_sc_hd__and2b_1 _14137_ (.A_N(_06872_),
    .B(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__a21o_1 _14138_ (.A1(_06860_),
    .A2(_06874_),
    .B1(_06872_),
    .X(_06875_));
 sky130_fd_sc_hd__xnor2_1 _14139_ (.A(_06859_),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__or2b_1 _14140_ (.A(_06859_),
    .B_N(_06875_),
    .X(_06877_));
 sky130_fd_sc_hd__a21boi_1 _14141_ (.A1(_06858_),
    .A2(_06876_),
    .B1_N(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__xor2_1 _14142_ (.A(_06857_),
    .B(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__nor2_1 _14143_ (.A(_06857_),
    .B(_06878_),
    .Y(_06880_));
 sky130_fd_sc_hd__a21oi_2 _14144_ (.A1(_06856_),
    .A2(_06879_),
    .B1(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_2 _14145_ (.A(_06842_),
    .B(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__and2_1 _14146_ (.A(_06842_),
    .B(_06881_),
    .X(_06883_));
 sky130_fd_sc_hd__xnor2_1 _14147_ (.A(_06856_),
    .B(_06879_),
    .Y(_06884_));
 sky130_fd_sc_hd__xnor2_1 _14148_ (.A(_06858_),
    .B(_06876_),
    .Y(_06885_));
 sky130_fd_sc_hd__xnor2_1 _14149_ (.A(_06860_),
    .B(_06874_),
    .Y(_06886_));
 sky130_fd_sc_hd__xnor2_2 _14150_ (.A(_06862_),
    .B(_06869_),
    .Y(_06887_));
 sky130_fd_sc_hd__nor2_1 _14151_ (.A(_05825_),
    .B(_06678_),
    .Y(_06888_));
 sky130_fd_sc_hd__o22ai_1 _14152_ (.A1(_05825_),
    .A2(_06740_),
    .B1(_06678_),
    .B2(_06704_),
    .Y(_06889_));
 sky130_fd_sc_hd__a21bo_1 _14153_ (.A1(_06741_),
    .A2(_06888_),
    .B1_N(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__nor2_1 _14154_ (.A(_06666_),
    .B(_06672_),
    .Y(_06891_));
 sky130_fd_sc_hd__xnor2_1 _14155_ (.A(_06890_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__xnor2_1 _14156_ (.A(_06865_),
    .B(_06867_),
    .Y(_06893_));
 sky130_fd_sc_hd__nor2_1 _14157_ (.A(_06805_),
    .B(_06663_),
    .Y(_06894_));
 sky130_fd_sc_hd__nor2_1 _14158_ (.A(_06776_),
    .B(_06677_),
    .Y(_06895_));
 sky130_fd_sc_hd__xor2_1 _14159_ (.A(_06864_),
    .B(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__and2_1 _14160_ (.A(_06864_),
    .B(_06895_),
    .X(_06897_));
 sky130_fd_sc_hd__a21oi_1 _14161_ (.A1(_06894_),
    .A2(_06896_),
    .B1(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__nand2_1 _14162_ (.A(_06893_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__nor2_1 _14163_ (.A(_06893_),
    .B(_06898_),
    .Y(_06900_));
 sky130_fd_sc_hd__a21oi_1 _14164_ (.A1(_06892_),
    .A2(_06899_),
    .B1(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__o22a_1 _14165_ (.A1(_06680_),
    .A2(_06690_),
    .B1(_06672_),
    .B2(_06675_),
    .X(_06902_));
 sky130_fd_sc_hd__or2_1 _14166_ (.A(_06853_),
    .B(_06902_),
    .X(_06903_));
 sky130_fd_sc_hd__a22o_1 _14167_ (.A1(_06741_),
    .A2(_06888_),
    .B1(_06889_),
    .B2(_06891_),
    .X(_06904_));
 sky130_fd_sc_hd__and2b_1 _14168_ (.A_N(_06903_),
    .B(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__and2b_1 _14169_ (.A_N(_06904_),
    .B(_06903_),
    .X(_06906_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(_06905_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__xor2_1 _14171_ (.A(_06887_),
    .B(_06901_),
    .X(_06908_));
 sky130_fd_sc_hd__nand2_1 _14172_ (.A(_06907_),
    .B(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__o21a_1 _14173_ (.A1(_06887_),
    .A2(_06901_),
    .B1(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__or2_1 _14174_ (.A(_06886_),
    .B(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__nand2_1 _14175_ (.A(_06886_),
    .B(_06910_),
    .Y(_06912_));
 sky130_fd_sc_hd__and2_1 _14176_ (.A(_06911_),
    .B(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__nand2_1 _14177_ (.A(_06905_),
    .B(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__and3_1 _14178_ (.A(_06885_),
    .B(_06911_),
    .C(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__or2_1 _14179_ (.A(_06905_),
    .B(_06913_),
    .X(_06916_));
 sky130_fd_sc_hd__nand2_1 _14180_ (.A(_06914_),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__nor2_1 _14181_ (.A(_06704_),
    .B(_06672_),
    .Y(_06918_));
 sky130_fd_sc_hd__nand2_1 _14182_ (.A(_06709_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__or2_1 _14183_ (.A(_06709_),
    .B(_06918_),
    .X(_06920_));
 sky130_fd_sc_hd__nand2_1 _14184_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__nor2_1 _14185_ (.A(_06666_),
    .B(_06690_),
    .Y(_06922_));
 sky130_fd_sc_hd__xnor2_1 _14186_ (.A(_06921_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__xnor2_1 _14187_ (.A(_06894_),
    .B(_06896_),
    .Y(_06924_));
 sky130_fd_sc_hd__nor2_1 _14188_ (.A(_06769_),
    .B(_06671_),
    .Y(_06925_));
 sky130_fd_sc_hd__nor2_1 _14189_ (.A(_05984_),
    .B(_06671_),
    .Y(_06926_));
 sky130_fd_sc_hd__o21ba_1 _14190_ (.A1(_06769_),
    .A2(_06677_),
    .B1_N(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__a21oi_1 _14191_ (.A1(_06895_),
    .A2(_06925_),
    .B1(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__or3b_1 _14192_ (.A(_06805_),
    .B(_06667_),
    .C_N(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__a21bo_1 _14193_ (.A1(_06895_),
    .A2(_06925_),
    .B1_N(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__xnor2_1 _14194_ (.A(_06924_),
    .B(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__xnor2_1 _14195_ (.A(_06923_),
    .B(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__o21bai_1 _14196_ (.A1(_06805_),
    .A2(_06668_),
    .B1_N(_06928_),
    .Y(_06933_));
 sky130_fd_sc_hd__nand2_1 _14197_ (.A(_06929_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__nor2_1 _14198_ (.A(_06769_),
    .B(_06610_),
    .Y(_06935_));
 sky130_fd_sc_hd__o22a_1 _14199_ (.A1(_06776_),
    .A2(_06610_),
    .B1(_06671_),
    .B2(_06769_),
    .X(_06936_));
 sky130_fd_sc_hd__a21oi_1 _14200_ (.A1(_06926_),
    .A2(_06935_),
    .B1(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__or3b_1 _14201_ (.A(_06805_),
    .B(_06678_),
    .C_N(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__a21boi_1 _14202_ (.A1(_06926_),
    .A2(_06935_),
    .B1_N(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__nor2_1 _14203_ (.A(_05825_),
    .B(_06690_),
    .Y(_06940_));
 sky130_fd_sc_hd__o22a_1 _14204_ (.A1(_06704_),
    .A2(_06690_),
    .B1(_06663_),
    .B2(_05825_),
    .X(_06941_));
 sky130_fd_sc_hd__a21oi_1 _14205_ (.A1(_06664_),
    .A2(_06940_),
    .B1(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__xor2_1 _14206_ (.A(_06934_),
    .B(_06939_),
    .X(_06943_));
 sky130_fd_sc_hd__nand2_1 _14207_ (.A(_06942_),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__o21ai_1 _14208_ (.A1(_06934_),
    .A2(_06939_),
    .B1(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__or2b_1 _14209_ (.A(_06932_),
    .B_N(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__nand2_1 _14210_ (.A(_06664_),
    .B(_06940_),
    .Y(_06947_));
 sky130_fd_sc_hd__xnor2_1 _14211_ (.A(_06932_),
    .B(_06945_),
    .Y(_06948_));
 sky130_fd_sc_hd__or2b_1 _14212_ (.A(_06947_),
    .B_N(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__o31a_1 _14213_ (.A1(_06666_),
    .A2(_06690_),
    .A3(_06921_),
    .B1(_06919_),
    .X(_06950_));
 sky130_fd_sc_hd__and2b_1 _14214_ (.A_N(_06950_),
    .B(_06852_),
    .X(_06951_));
 sky130_fd_sc_hd__and2b_1 _14215_ (.A_N(_06852_),
    .B(_06950_),
    .X(_06952_));
 sky130_fd_sc_hd__nor2_1 _14216_ (.A(_06951_),
    .B(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__and2b_1 _14217_ (.A_N(_06900_),
    .B(_06899_),
    .X(_06954_));
 sky130_fd_sc_hd__xnor2_1 _14218_ (.A(_06892_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__or2b_1 _14219_ (.A(_06924_),
    .B_N(_06930_),
    .X(_06956_));
 sky130_fd_sc_hd__a21boi_1 _14220_ (.A1(_06923_),
    .A2(_06931_),
    .B1_N(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__nor2_1 _14221_ (.A(_06955_),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__nand2_1 _14222_ (.A(_06955_),
    .B(_06957_),
    .Y(_06959_));
 sky130_fd_sc_hd__and2b_1 _14223_ (.A_N(_06958_),
    .B(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__xnor2_1 _14224_ (.A(_06953_),
    .B(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__a21oi_1 _14225_ (.A1(_06946_),
    .A2(_06949_),
    .B1(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__nor2_1 _14226_ (.A(_06805_),
    .B(_06672_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand2_1 _14227_ (.A(_06935_),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__or2_1 _14228_ (.A(_06935_),
    .B(_06963_),
    .X(_06965_));
 sky130_fd_sc_hd__and2_1 _14229_ (.A(_06964_),
    .B(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__nand2_1 _14230_ (.A(_06888_),
    .B(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__o211ai_1 _14231_ (.A1(_06888_),
    .A2(_06966_),
    .B1(_06963_),
    .C1(_06940_),
    .Y(_06968_));
 sky130_fd_sc_hd__or2_1 _14232_ (.A(_06942_),
    .B(_06943_),
    .X(_06969_));
 sky130_fd_sc_hd__nand2_1 _14233_ (.A(_06944_),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__o21bai_1 _14234_ (.A1(_06805_),
    .A2(_06678_),
    .B1_N(_06937_),
    .Y(_06971_));
 sky130_fd_sc_hd__and2_1 _14235_ (.A(_06938_),
    .B(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__xnor2_1 _14236_ (.A(_06964_),
    .B(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__and2_1 _14237_ (.A(_06844_),
    .B(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__a31o_1 _14238_ (.A1(_06935_),
    .A2(_06963_),
    .A3(_06972_),
    .B1(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__xor2_1 _14239_ (.A(_06970_),
    .B(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__nor2_1 _14240_ (.A(_06844_),
    .B(_06973_),
    .Y(_06977_));
 sky130_fd_sc_hd__or2_1 _14241_ (.A(_06974_),
    .B(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__a211oi_1 _14242_ (.A1(_06967_),
    .A2(_06968_),
    .B1(_06976_),
    .C1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__xor2_1 _14243_ (.A(_06947_),
    .B(_06948_),
    .X(_06980_));
 sky130_fd_sc_hd__a21oi_1 _14244_ (.A1(_06946_),
    .A2(_06961_),
    .B1(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__and3b_1 _14245_ (.A_N(_06962_),
    .B(_06979_),
    .C(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__and3_1 _14246_ (.A(_06944_),
    .B(_06969_),
    .C(_06975_),
    .X(_06983_));
 sky130_fd_sc_hd__and2_1 _14247_ (.A(_06981_),
    .B(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__or2_1 _14248_ (.A(_06907_),
    .B(_06908_),
    .X(_06985_));
 sky130_fd_sc_hd__nand2_1 _14249_ (.A(_06909_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__a21o_1 _14250_ (.A1(_06953_),
    .A2(_06959_),
    .B1(_06958_),
    .X(_06987_));
 sky130_fd_sc_hd__xnor2_1 _14251_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__or4_1 _14252_ (.A(_06951_),
    .B(_06962_),
    .C(_06984_),
    .D(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__and2b_1 _14253_ (.A_N(_06986_),
    .B(_06987_),
    .X(_06990_));
 sky130_fd_sc_hd__a21o_1 _14254_ (.A1(_06951_),
    .A2(_06988_),
    .B1(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__o22a_1 _14255_ (.A1(_06962_),
    .A2(_06984_),
    .B1(_06988_),
    .B2(_06951_),
    .X(_06992_));
 sky130_fd_sc_hd__a211oi_1 _14256_ (.A1(_06982_),
    .A2(_06989_),
    .B1(_06991_),
    .C1(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__or4_2 _14257_ (.A(_06884_),
    .B(_06915_),
    .C(_06917_),
    .D(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__nor3_4 _14258_ (.A(_06882_),
    .B(_06883_),
    .C(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nor2_1 _14259_ (.A(_06724_),
    .B(_06672_),
    .Y(_06996_));
 sky130_fd_sc_hd__or2_1 _14260_ (.A(_06134_),
    .B(_06667_),
    .X(_06997_));
 sky130_fd_sc_hd__xnor2_1 _14261_ (.A(_06997_),
    .B(_06725_),
    .Y(_06998_));
 sky130_fd_sc_hd__xnor2_1 _14262_ (.A(_06996_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__o31a_1 _14263_ (.A1(_06698_),
    .A2(_06726_),
    .A3(_06672_),
    .B1(_06729_),
    .X(_07000_));
 sky130_fd_sc_hd__nor2_1 _14264_ (.A(_06999_),
    .B(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__and2_1 _14265_ (.A(_06999_),
    .B(_07000_),
    .X(_07002_));
 sky130_fd_sc_hd__or2_2 _14266_ (.A(_07001_),
    .B(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__a21oi_2 _14267_ (.A1(_06744_),
    .A2(_06751_),
    .B1(_06755_),
    .Y(_07004_));
 sky130_fd_sc_hd__xnor2_2 _14268_ (.A(_07003_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__xnor2_2 _14269_ (.A(_07005_),
    .B(_06732_),
    .Y(_07006_));
 sky130_fd_sc_hd__a21bo_1 _14270_ (.A1(_06762_),
    .A2(_06765_),
    .B1_N(_06764_),
    .X(_07007_));
 sky130_fd_sc_hd__nor2_1 _14271_ (.A(_06245_),
    .B(_06663_),
    .Y(_07008_));
 sky130_fd_sc_hd__nor2_1 _14272_ (.A(_06675_),
    .B(_06740_),
    .Y(_07009_));
 sky130_fd_sc_hd__nor2_1 _14273_ (.A(_06680_),
    .B(_06708_),
    .Y(_07010_));
 sky130_fd_sc_hd__xnor2_1 _14274_ (.A(_07009_),
    .B(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__xnor2_1 _14275_ (.A(_07008_),
    .B(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__xnor2_2 _14276_ (.A(_07007_),
    .B(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__o31a_1 _14277_ (.A1(_06689_),
    .A2(_06668_),
    .A3(_06750_),
    .B1(_06748_),
    .X(_07014_));
 sky130_fd_sc_hd__xor2_2 _14278_ (.A(_07013_),
    .B(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__nor2_1 _14279_ (.A(_06666_),
    .B(_06760_),
    .Y(_07016_));
 sky130_fd_sc_hd__xnor2_2 _14280_ (.A(_06705_),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__o21ai_1 _14281_ (.A1(_06805_),
    .A2(_06761_),
    .B1(_06772_),
    .Y(_07018_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(_06774_),
    .B(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__xor2_2 _14283_ (.A(_07017_),
    .B(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__a31o_1 _14284_ (.A1(_06766_),
    .A2(_06767_),
    .A3(_06782_),
    .B1(_06781_),
    .X(_07021_));
 sky130_fd_sc_hd__xor2_2 _14285_ (.A(_07020_),
    .B(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__xnor2_2 _14286_ (.A(_07015_),
    .B(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__or2b_1 _14287_ (.A(_06784_),
    .B_N(_06796_),
    .X(_07024_));
 sky130_fd_sc_hd__a21boi_2 _14288_ (.A1(_06757_),
    .A2(_06797_),
    .B1_N(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__xor2_2 _14289_ (.A(_07023_),
    .B(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__xnor2_2 _14290_ (.A(_07006_),
    .B(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__or2b_1 _14291_ (.A(_06798_),
    .B_N(_06816_),
    .X(_07028_));
 sky130_fd_sc_hd__a21boi_2 _14292_ (.A1(_06737_),
    .A2(_06817_),
    .B1_N(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__xor2_2 _14293_ (.A(_07027_),
    .B(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__xnor2_2 _14294_ (.A(_06735_),
    .B(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__nor2_1 _14295_ (.A(_06818_),
    .B(_06840_),
    .Y(_07032_));
 sky130_fd_sc_hd__a21oi_2 _14296_ (.A1(_06703_),
    .A2(_06841_),
    .B1(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__xor2_2 _14297_ (.A(_07031_),
    .B(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__and2_1 _14298_ (.A(_06882_),
    .B(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__xor2_1 _14299_ (.A(_06842_),
    .B(_06881_),
    .X(_07036_));
 sky130_fd_sc_hd__a211oi_2 _14300_ (.A1(_06911_),
    .A2(_06914_),
    .B1(_06884_),
    .C1(_06885_),
    .Y(_07037_));
 sky130_fd_sc_hd__and3_1 _14301_ (.A(_07034_),
    .B(_07036_),
    .C(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__a211o_1 _14302_ (.A1(_07036_),
    .A2(_07037_),
    .B1(_06882_),
    .C1(_07034_),
    .X(_07039_));
 sky130_fd_sc_hd__nor3b_2 _14303_ (.A(_07035_),
    .B(_07038_),
    .C_N(_07039_),
    .Y(_07040_));
 sky130_fd_sc_hd__xor2_4 _14304_ (.A(_06995_),
    .B(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__nand2_1 _14305_ (.A(_06882_),
    .B(_07034_),
    .Y(_07042_));
 sky130_fd_sc_hd__a31o_1 _14306_ (.A1(_07042_),
    .A2(_06995_),
    .A3(_07039_),
    .B1(_07038_),
    .X(_07043_));
 sky130_fd_sc_hd__o32ai_4 _14307_ (.A1(_07005_),
    .A2(_06731_),
    .A3(_06700_),
    .B1(_07004_),
    .B2(_07003_),
    .Y(_07044_));
 sky130_fd_sc_hd__nor2_1 _14308_ (.A(_06134_),
    .B(_06662_),
    .Y(_07045_));
 sky130_fd_sc_hd__nor2_1 _14309_ (.A(_06696_),
    .B(_06667_),
    .Y(_07046_));
 sky130_fd_sc_hd__xor2_1 _14310_ (.A(_07045_),
    .B(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__or3b_1 _14311_ (.A(_06067_),
    .B(_06678_),
    .C_N(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__o21bai_1 _14312_ (.A1(_06724_),
    .A2(_06678_),
    .B1_N(_07047_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand2_1 _14313_ (.A(_07048_),
    .B(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__nand2_1 _14314_ (.A(_06996_),
    .B(_06998_),
    .Y(_07051_));
 sky130_fd_sc_hd__o21a_1 _14315_ (.A1(_06997_),
    .A2(_06726_),
    .B1(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__nor2_1 _14316_ (.A(_07050_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__and2_1 _14317_ (.A(_07050_),
    .B(_07052_),
    .X(_07054_));
 sky130_fd_sc_hd__or2_1 _14318_ (.A(_07053_),
    .B(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__nand2_1 _14319_ (.A(_07007_),
    .B(_07012_),
    .Y(_07056_));
 sky130_fd_sc_hd__o21a_1 _14320_ (.A1(_07013_),
    .A2(_07014_),
    .B1(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__xnor2_1 _14321_ (.A(_07055_),
    .B(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__xnor2_1 _14322_ (.A(_07058_),
    .B(_07001_),
    .Y(_07059_));
 sky130_fd_sc_hd__nor2_1 _14323_ (.A(_05982_),
    .B(_06658_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_1 _14324_ (.A(_07060_),
    .B(_06843_),
    .Y(_07061_));
 sky130_fd_sc_hd__or2_1 _14325_ (.A(_06245_),
    .B(_06708_),
    .X(_07062_));
 sky130_fd_sc_hd__and3b_1 _14326_ (.A_N(_06240_),
    .B(_06758_),
    .C(_06759_),
    .X(_07063_));
 sky130_fd_sc_hd__or2_1 _14327_ (.A(_06680_),
    .B(_06739_),
    .X(_07064_));
 sky130_fd_sc_hd__xnor2_1 _14328_ (.A(_07063_),
    .B(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__xnor2_1 _14329_ (.A(_07062_),
    .B(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__xor2_1 _14330_ (.A(_07061_),
    .B(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__or3_1 _14331_ (.A(_06689_),
    .B(_06663_),
    .C(_07011_),
    .X(_07068_));
 sky130_fd_sc_hd__o31a_1 _14332_ (.A1(_06675_),
    .A2(_06708_),
    .A3(_07064_),
    .B1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__xor2_1 _14333_ (.A(_07067_),
    .B(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__xor2_1 _14334_ (.A(_06705_),
    .B(_07060_),
    .X(_07071_));
 sky130_fd_sc_hd__buf_2 _14335_ (.A(_06658_),
    .X(_07072_));
 sky130_fd_sc_hd__or2_1 _14336_ (.A(_06776_),
    .B(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__a21oi_1 _14337_ (.A1(_06017_),
    .A2(_07073_),
    .B1(_06770_),
    .Y(_07074_));
 sky130_fd_sc_hd__nand2_1 _14338_ (.A(_07071_),
    .B(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__or2_1 _14339_ (.A(_07071_),
    .B(_07074_),
    .X(_07076_));
 sky130_fd_sc_hd__and2_1 _14340_ (.A(_07075_),
    .B(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__o21ai_1 _14341_ (.A1(_07017_),
    .A2(_07019_),
    .B1(_06774_),
    .Y(_07078_));
 sky130_fd_sc_hd__xor2_1 _14342_ (.A(_07077_),
    .B(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__xnor2_1 _14343_ (.A(_07070_),
    .B(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__and2_1 _14344_ (.A(_07020_),
    .B(_07021_),
    .X(_07081_));
 sky130_fd_sc_hd__a21oi_1 _14345_ (.A1(_07015_),
    .A2(_07022_),
    .B1(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__xor2_1 _14346_ (.A(_07080_),
    .B(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__nand2_1 _14347_ (.A(_07059_),
    .B(_07083_),
    .Y(_07084_));
 sky130_fd_sc_hd__or2_1 _14348_ (.A(_07059_),
    .B(_07083_),
    .X(_07085_));
 sky130_fd_sc_hd__nand2_1 _14349_ (.A(_07084_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__nor2_1 _14350_ (.A(_07023_),
    .B(_07025_),
    .Y(_07087_));
 sky130_fd_sc_hd__a21oi_1 _14351_ (.A1(_07006_),
    .A2(_07026_),
    .B1(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__xor2_1 _14352_ (.A(_07086_),
    .B(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__xnor2_1 _14353_ (.A(_07044_),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__nor2_1 _14354_ (.A(_07027_),
    .B(_07029_),
    .Y(_07091_));
 sky130_fd_sc_hd__a21oi_1 _14355_ (.A1(_06735_),
    .A2(_07030_),
    .B1(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__nor2_1 _14356_ (.A(_07090_),
    .B(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__and2_1 _14357_ (.A(_07090_),
    .B(_07092_),
    .X(_07094_));
 sky130_fd_sc_hd__nor2_2 _14358_ (.A(_07093_),
    .B(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__nor2_1 _14359_ (.A(_07031_),
    .B(_07033_),
    .Y(_07096_));
 sky130_fd_sc_hd__a21oi_1 _14360_ (.A1(_06882_),
    .A2(_07034_),
    .B1(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__xnor2_1 _14361_ (.A(_07095_),
    .B(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__and2_1 _14362_ (.A(_07043_),
    .B(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__nor2_1 _14363_ (.A(_07043_),
    .B(_07098_),
    .Y(_07100_));
 sky130_fd_sc_hd__or2_1 _14364_ (.A(_07099_),
    .B(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__nor2_1 _14365_ (.A(_05793_),
    .B(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__a21oi_1 _14366_ (.A1(_05793_),
    .A2(_07041_),
    .B1(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__or2_2 _14367_ (.A(_05779_),
    .B(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__inv_2 _14368_ (.A(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__buf_2 _14369_ (.A(_05931_),
    .X(_07106_));
 sky130_fd_sc_hd__clkbuf_4 _14370_ (.A(_05893_),
    .X(_07107_));
 sky130_fd_sc_hd__or2_2 _14371_ (.A(_06680_),
    .B(_07072_),
    .X(_07108_));
 sky130_fd_sc_hd__or2_1 _14372_ (.A(_06240_),
    .B(_06658_),
    .X(_07109_));
 sky130_fd_sc_hd__xnor2_2 _14373_ (.A(_07108_),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__nor2_1 _14374_ (.A(_06689_),
    .B(_07072_),
    .Y(_07111_));
 sky130_fd_sc_hd__xor2_1 _14375_ (.A(_07110_),
    .B(_07111_),
    .X(_07112_));
 sky130_fd_sc_hd__o32a_1 _14376_ (.A1(_06689_),
    .A2(_06760_),
    .A3(_07110_),
    .B1(_07108_),
    .B2(_06675_),
    .X(_07113_));
 sky130_fd_sc_hd__nor2_1 _14377_ (.A(_07112_),
    .B(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__or2_1 _14378_ (.A(_06724_),
    .B(_06740_),
    .X(_07115_));
 sky130_fd_sc_hd__nor2_1 _14379_ (.A(_06698_),
    .B(_07072_),
    .Y(_07116_));
 sky130_fd_sc_hd__and2_1 _14380_ (.A(_06176_),
    .B(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__o21ba_1 _14381_ (.A1(_06696_),
    .A2(_06760_),
    .B1_N(_07116_),
    .X(_07118_));
 sky130_fd_sc_hd__or2_1 _14382_ (.A(_07117_),
    .B(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__xnor2_1 _14383_ (.A(_07115_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__or2_1 _14384_ (.A(_06696_),
    .B(_06740_),
    .X(_07121_));
 sky130_fd_sc_hd__or2_1 _14385_ (.A(_06724_),
    .B(_06708_),
    .X(_07122_));
 sky130_fd_sc_hd__nor2_1 _14386_ (.A(_06698_),
    .B(_06760_),
    .Y(_07123_));
 sky130_fd_sc_hd__xnor2_1 _14387_ (.A(_07121_),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__or2b_1 _14388_ (.A(_07122_),
    .B_N(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__o31a_1 _14389_ (.A1(_06698_),
    .A2(_07121_),
    .A3(_06760_),
    .B1(_07125_),
    .X(_07126_));
 sky130_fd_sc_hd__xor2_1 _14390_ (.A(_07120_),
    .B(_07126_),
    .X(_07127_));
 sky130_fd_sc_hd__o21ai_1 _14391_ (.A1(_06675_),
    .A2(_06761_),
    .B1(_07108_),
    .Y(_07128_));
 sky130_fd_sc_hd__or2_1 _14392_ (.A(_07111_),
    .B(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__o32ai_1 _14393_ (.A1(_06689_),
    .A2(_07072_),
    .A3(_07110_),
    .B1(_07108_),
    .B2(_06675_),
    .Y(_07130_));
 sky130_fd_sc_hd__nand2_1 _14394_ (.A(_07111_),
    .B(_07128_),
    .Y(_07131_));
 sky130_fd_sc_hd__nand2_1 _14395_ (.A(_07130_),
    .B(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__a21oi_1 _14396_ (.A1(_07129_),
    .A2(_07132_),
    .B1(_06239_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_1 _14397_ (.A(_07114_),
    .B(_07127_),
    .Y(_07134_));
 sky130_fd_sc_hd__or2_1 _14398_ (.A(_07114_),
    .B(_07127_),
    .X(_07135_));
 sky130_fd_sc_hd__nor2_1 _14399_ (.A(_06698_),
    .B(_06740_),
    .Y(_07136_));
 sky130_fd_sc_hd__nor2_1 _14400_ (.A(_06696_),
    .B(_06708_),
    .Y(_07137_));
 sky130_fd_sc_hd__xnor2_1 _14401_ (.A(_07136_),
    .B(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__nor3_1 _14402_ (.A(_06724_),
    .B(_06663_),
    .C(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__a21oi_1 _14403_ (.A1(_07136_),
    .A2(_07137_),
    .B1(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__xnor2_1 _14404_ (.A(_07122_),
    .B(_07124_),
    .Y(_07141_));
 sky130_fd_sc_hd__and2b_1 _14405_ (.A_N(_07140_),
    .B(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__a21oi_1 _14406_ (.A1(_07134_),
    .A2(_07135_),
    .B1(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__or2_1 _14407_ (.A(_07133_),
    .B(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__nor2_1 _14408_ (.A(_06680_),
    .B(_06761_),
    .Y(_07145_));
 sky130_fd_sc_hd__o31a_1 _14409_ (.A1(_06239_),
    .A2(_07111_),
    .A3(_07145_),
    .B1(_07131_),
    .X(_07146_));
 sky130_fd_sc_hd__or2_1 _14410_ (.A(_07120_),
    .B(_07126_),
    .X(_07147_));
 sky130_fd_sc_hd__o21ba_1 _14411_ (.A1(_07115_),
    .A2(_07119_),
    .B1_N(_07117_),
    .X(_07148_));
 sky130_fd_sc_hd__a21oi_1 _14412_ (.A1(_06696_),
    .A2(_06698_),
    .B1(_07072_),
    .Y(_07149_));
 sky130_fd_sc_hd__or3b_1 _14413_ (.A(_06760_),
    .B(_07117_),
    .C_N(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__and3b_1 _14414_ (.A_N(_07072_),
    .B(_07148_),
    .C(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__xnor2_1 _14415_ (.A(_07132_),
    .B(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__xnor2_1 _14416_ (.A(_07147_),
    .B(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__and2_1 _14417_ (.A(_07146_),
    .B(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__nor2_1 _14418_ (.A(_07146_),
    .B(_07153_),
    .Y(_07155_));
 sky130_fd_sc_hd__or2_1 _14419_ (.A(_07154_),
    .B(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__xor2_1 _14420_ (.A(_07144_),
    .B(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__and3_1 _14421_ (.A(_07114_),
    .B(_07127_),
    .C(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__a21oi_1 _14422_ (.A1(_07114_),
    .A2(_07127_),
    .B1(_07157_),
    .Y(_07159_));
 sky130_fd_sc_hd__or2_1 _14423_ (.A(_07158_),
    .B(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__nand2_1 _14424_ (.A(_07133_),
    .B(_07143_),
    .Y(_07161_));
 sky130_fd_sc_hd__nand2_1 _14425_ (.A(_07144_),
    .B(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__o21a_1 _14426_ (.A1(_06724_),
    .A2(_06663_),
    .B1(_07138_),
    .X(_07163_));
 sky130_fd_sc_hd__or2_1 _14427_ (.A(_07139_),
    .B(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__or2_1 _14428_ (.A(_06067_),
    .B(_06668_),
    .X(_07165_));
 sky130_fd_sc_hd__o22a_1 _14429_ (.A1(_06696_),
    .A2(_06663_),
    .B1(_06708_),
    .B2(_06698_),
    .X(_07166_));
 sky130_fd_sc_hd__o2bb2a_1 _14430_ (.A1_N(_07137_),
    .A2_N(_07045_),
    .B1(_07165_),
    .B2(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__or2_1 _14431_ (.A(_07164_),
    .B(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__and2b_1 _14432_ (.A_N(_07141_),
    .B(_07140_),
    .X(_07169_));
 sky130_fd_sc_hd__or2_1 _14433_ (.A(_07142_),
    .B(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__and2_1 _14434_ (.A(_06153_),
    .B(_06705_),
    .X(_07171_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14435_ (.A(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__nor2_1 _14436_ (.A(_06689_),
    .B(_06760_),
    .Y(_07173_));
 sky130_fd_sc_hd__xnor2_1 _14437_ (.A(_07110_),
    .B(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__xnor2_1 _14438_ (.A(_07172_),
    .B(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__nor2_1 _14439_ (.A(_06689_),
    .B(_06740_),
    .Y(_07176_));
 sky130_fd_sc_hd__and3b_1 _14440_ (.A_N(_06680_),
    .B(_06758_),
    .C(_06759_),
    .X(_07177_));
 sky130_fd_sc_hd__xnor2_1 _14441_ (.A(_07109_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__and2b_1 _14442_ (.A_N(_07108_),
    .B(_07063_),
    .X(_07179_));
 sky130_fd_sc_hd__a21oi_1 _14443_ (.A1(_07176_),
    .A2(_07178_),
    .B1(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_1 _14444_ (.A(_07172_),
    .B(_07174_),
    .Y(_07181_));
 sky130_fd_sc_hd__o21a_1 _14445_ (.A1(_07175_),
    .A2(_07180_),
    .B1(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__xor2_1 _14446_ (.A(_07170_),
    .B(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__xnor2_1 _14447_ (.A(_07168_),
    .B(_07183_),
    .Y(_07184_));
 sky130_fd_sc_hd__and2_1 _14448_ (.A(_07112_),
    .B(_07113_),
    .X(_07185_));
 sky130_fd_sc_hd__nor2_1 _14449_ (.A(_07114_),
    .B(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__a21o_1 _14450_ (.A1(_06153_),
    .A2(_07072_),
    .B1(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__o21ba_1 _14451_ (.A1(_06704_),
    .A2(_06761_),
    .B1_N(_07060_),
    .X(_07188_));
 sky130_fd_sc_hd__xor2_1 _14452_ (.A(_07175_),
    .B(_07180_),
    .X(_07189_));
 sky130_fd_sc_hd__and2b_1 _14453_ (.A_N(_07188_),
    .B(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__and2_1 _14454_ (.A(_07187_),
    .B(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__nor2_1 _14455_ (.A(_07187_),
    .B(_07190_),
    .Y(_07192_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_07191_),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__a21oi_1 _14457_ (.A1(_07184_),
    .A2(_07193_),
    .B1(_07191_),
    .Y(_07194_));
 sky130_fd_sc_hd__xnor2_1 _14458_ (.A(_07162_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__or2b_1 _14459_ (.A(_07168_),
    .B_N(_07183_),
    .X(_07196_));
 sky130_fd_sc_hd__o21ai_1 _14460_ (.A1(_07170_),
    .A2(_07182_),
    .B1(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__or2b_1 _14461_ (.A(_07195_),
    .B_N(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__o21a_1 _14462_ (.A1(_07162_),
    .A2(_07194_),
    .B1(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__nor2_1 _14463_ (.A(_07160_),
    .B(_07199_),
    .Y(_07200_));
 sky130_fd_sc_hd__inv_2 _14464_ (.A(_07151_),
    .Y(_07201_));
 sky130_fd_sc_hd__or2b_1 _14465_ (.A(_07147_),
    .B_N(_07152_),
    .X(_07202_));
 sky130_fd_sc_hd__o21ai_1 _14466_ (.A1(_07132_),
    .A2(_07201_),
    .B1(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__or2_1 _14467_ (.A(_06689_),
    .B(_06761_),
    .X(_07204_));
 sky130_fd_sc_hd__or3_1 _14468_ (.A(_06724_),
    .B(_06760_),
    .C(_07117_),
    .X(_07205_));
 sky130_fd_sc_hd__nor2_1 _14469_ (.A(_07131_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__and2_1 _14470_ (.A(_07131_),
    .B(_07205_),
    .X(_07207_));
 sky130_fd_sc_hd__or2_1 _14471_ (.A(_07206_),
    .B(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__xnor2_1 _14472_ (.A(_07148_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__a21oi_1 _14473_ (.A1(_07204_),
    .A2(_07209_),
    .B1(_07154_),
    .Y(_07210_));
 sky130_fd_sc_hd__xnor2_1 _14474_ (.A(_07203_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ba_1 _14475_ (.A1(_07144_),
    .A2(_07156_),
    .B1_N(_07158_),
    .X(_07212_));
 sky130_fd_sc_hd__nor2_1 _14476_ (.A(_07211_),
    .B(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__and2_1 _14477_ (.A(_07211_),
    .B(_07212_),
    .X(_07214_));
 sky130_fd_sc_hd__nor2_1 _14478_ (.A(_07213_),
    .B(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__and2_1 _14479_ (.A(_07200_),
    .B(_07215_),
    .X(_07216_));
 sky130_fd_sc_hd__nor2_1 _14480_ (.A(_07200_),
    .B(_07215_),
    .Y(_07217_));
 sky130_fd_sc_hd__nor2_2 _14481_ (.A(_07216_),
    .B(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__nand2_1 _14482_ (.A(_07164_),
    .B(_07167_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_1 _14483_ (.A(_07168_),
    .B(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__xor2_1 _14484_ (.A(_07176_),
    .B(_07178_),
    .X(_07221_));
 sky130_fd_sc_hd__xnor2_1 _14485_ (.A(_07172_),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__nor2_1 _14486_ (.A(_06689_),
    .B(_06708_),
    .Y(_07223_));
 sky130_fd_sc_hd__a22o_1 _14487_ (.A1(_07177_),
    .A2(_07009_),
    .B1(_07223_),
    .B2(_07065_),
    .X(_07224_));
 sky130_fd_sc_hd__and2b_1 _14488_ (.A_N(_07222_),
    .B(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__a21oi_1 _14489_ (.A1(_07172_),
    .A2(_07221_),
    .B1(_07225_),
    .Y(_07226_));
 sky130_fd_sc_hd__xor2_1 _14490_ (.A(_07220_),
    .B(_07226_),
    .X(_07227_));
 sky130_fd_sc_hd__a21o_1 _14491_ (.A1(_07137_),
    .A2(_07045_),
    .B1(_07166_),
    .X(_07228_));
 sky130_fd_sc_hd__xnor2_1 _14492_ (.A(_07165_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__a21bo_1 _14493_ (.A1(_07045_),
    .A2(_07046_),
    .B1_N(_07048_),
    .X(_07230_));
 sky130_fd_sc_hd__and2b_1 _14494_ (.A_N(_07229_),
    .B(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__nor2_1 _14495_ (.A(_07220_),
    .B(_07226_),
    .Y(_07232_));
 sky130_fd_sc_hd__a21o_1 _14496_ (.A1(_07227_),
    .A2(_07231_),
    .B1(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__xnor2_1 _14497_ (.A(_07184_),
    .B(_07193_),
    .Y(_07234_));
 sky130_fd_sc_hd__xor2_1 _14498_ (.A(_07227_),
    .B(_07231_),
    .X(_07235_));
 sky130_fd_sc_hd__xor2_1 _14499_ (.A(_07188_),
    .B(_07189_),
    .X(_07236_));
 sky130_fd_sc_hd__xnor2_1 _14500_ (.A(_07222_),
    .B(_07224_),
    .Y(_07237_));
 sky130_fd_sc_hd__nand2_1 _14501_ (.A(_06002_),
    .B(_07072_),
    .Y(_07238_));
 sky130_fd_sc_hd__nand2_1 _14502_ (.A(_06002_),
    .B(_06770_),
    .Y(_07239_));
 sky130_fd_sc_hd__or4bb_1 _14503_ (.A(_06239_),
    .B(_07071_),
    .C_N(_07238_),
    .D_N(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__nor2_1 _14504_ (.A(_06239_),
    .B(_07071_),
    .Y(_07241_));
 sky130_fd_sc_hd__a22o_1 _14505_ (.A1(_07238_),
    .A2(_07241_),
    .B1(_07239_),
    .B2(_07075_),
    .X(_07242_));
 sky130_fd_sc_hd__a21boi_1 _14506_ (.A1(_07237_),
    .A2(_07240_),
    .B1_N(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__nand2_1 _14507_ (.A(_07236_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__nor2_1 _14508_ (.A(_07236_),
    .B(_07243_),
    .Y(_07245_));
 sky130_fd_sc_hd__a21oi_1 _14509_ (.A1(_07235_),
    .A2(_07244_),
    .B1(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__nor2_1 _14510_ (.A(_07234_),
    .B(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__and2_1 _14511_ (.A(_07234_),
    .B(_07246_),
    .X(_07248_));
 sky130_fd_sc_hd__nor2_1 _14512_ (.A(_07247_),
    .B(_07248_),
    .Y(_07249_));
 sky130_fd_sc_hd__xnor2_1 _14513_ (.A(_07233_),
    .B(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__and2b_1 _14514_ (.A_N(_07245_),
    .B(_07244_),
    .X(_07251_));
 sky130_fd_sc_hd__xnor2_1 _14515_ (.A(_07235_),
    .B(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__nor2_1 _14516_ (.A(_07067_),
    .B(_07069_),
    .Y(_07253_));
 sky130_fd_sc_hd__a31o_1 _14517_ (.A1(_07060_),
    .A2(_06843_),
    .A3(_07066_),
    .B1(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__and2b_1 _14518_ (.A_N(_07230_),
    .B(_07229_),
    .X(_07255_));
 sky130_fd_sc_hd__o21a_1 _14519_ (.A1(_07231_),
    .A2(_07255_),
    .B1(_05752_),
    .X(_07256_));
 sky130_fd_sc_hd__inv_2 _14520_ (.A(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__xnor2_1 _14521_ (.A(_07254_),
    .B(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__xnor2_1 _14522_ (.A(_07258_),
    .B(_07053_),
    .Y(_07259_));
 sky130_fd_sc_hd__and2_1 _14523_ (.A(_07242_),
    .B(_07240_),
    .X(_07260_));
 sky130_fd_sc_hd__xnor2_1 _14524_ (.A(_07237_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__and2_1 _14525_ (.A(_07077_),
    .B(_07078_),
    .X(_07262_));
 sky130_fd_sc_hd__a21oi_1 _14526_ (.A1(_07070_),
    .A2(_07079_),
    .B1(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__nor2_1 _14527_ (.A(_07261_),
    .B(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__nand2_1 _14528_ (.A(_07261_),
    .B(_07263_),
    .Y(_07265_));
 sky130_fd_sc_hd__and2b_1 _14529_ (.A_N(_07264_),
    .B(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__a21oi_1 _14530_ (.A1(_07259_),
    .A2(_07266_),
    .B1(_07264_),
    .Y(_07267_));
 sky130_fd_sc_hd__xnor2_1 _14531_ (.A(_07252_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__nand2_1 _14532_ (.A(_07254_),
    .B(_07257_),
    .Y(_07269_));
 sky130_fd_sc_hd__o31ai_2 _14533_ (.A1(_07258_),
    .A2(_07050_),
    .A3(_07052_),
    .B1(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__or2b_1 _14534_ (.A(_07268_),
    .B_N(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__o21a_1 _14535_ (.A1(_07252_),
    .A2(_07267_),
    .B1(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__or2_1 _14536_ (.A(_07250_),
    .B(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__xor2_1 _14537_ (.A(_07197_),
    .B(_07195_),
    .X(_07274_));
 sky130_fd_sc_hd__a21oi_1 _14538_ (.A1(_07233_),
    .A2(_07249_),
    .B1(_07247_),
    .Y(_07275_));
 sky130_fd_sc_hd__nor2_1 _14539_ (.A(_07274_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__and2_1 _14540_ (.A(_07274_),
    .B(_07275_),
    .X(_07277_));
 sky130_fd_sc_hd__nor2_1 _14541_ (.A(_07276_),
    .B(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__or2b_1 _14542_ (.A(_07273_),
    .B_N(_07278_),
    .X(_07279_));
 sky130_fd_sc_hd__xor2_1 _14543_ (.A(_07160_),
    .B(_07199_),
    .X(_07280_));
 sky130_fd_sc_hd__and2_1 _14544_ (.A(_07276_),
    .B(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__nor2_1 _14545_ (.A(_07276_),
    .B(_07280_),
    .Y(_07282_));
 sky130_fd_sc_hd__nor2_1 _14546_ (.A(_07281_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__xnor2_1 _14547_ (.A(_07279_),
    .B(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__xor2_1 _14548_ (.A(_07250_),
    .B(_07272_),
    .X(_07285_));
 sky130_fd_sc_hd__xor2_1 _14549_ (.A(_07270_),
    .B(_07268_),
    .X(_07286_));
 sky130_fd_sc_hd__xnor2_1 _14550_ (.A(_07259_),
    .B(_07266_),
    .Y(_07287_));
 sky130_fd_sc_hd__o21a_1 _14551_ (.A1(_07080_),
    .A2(_07082_),
    .B1(_07084_),
    .X(_07288_));
 sky130_fd_sc_hd__o32ai_2 _14552_ (.A1(_07058_),
    .A2(_06999_),
    .A3(_07000_),
    .B1(_07057_),
    .B2(_07055_),
    .Y(_07289_));
 sky130_fd_sc_hd__xor2_1 _14553_ (.A(_07287_),
    .B(_07288_),
    .X(_07290_));
 sky130_fd_sc_hd__nand2_1 _14554_ (.A(_07289_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__o21a_1 _14555_ (.A1(_07287_),
    .A2(_07288_),
    .B1(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__nor2_1 _14556_ (.A(_07286_),
    .B(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__xor2_1 _14557_ (.A(_07285_),
    .B(_07293_),
    .X(_07294_));
 sky130_fd_sc_hd__xnor2_1 _14558_ (.A(_07286_),
    .B(_07292_),
    .Y(_07295_));
 sky130_fd_sc_hd__or2_1 _14559_ (.A(_07289_),
    .B(_07290_),
    .X(_07296_));
 sky130_fd_sc_hd__nand2_1 _14560_ (.A(_07291_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__nor2_1 _14561_ (.A(_07086_),
    .B(_07088_),
    .Y(_07298_));
 sky130_fd_sc_hd__a21oi_1 _14562_ (.A1(_07044_),
    .A2(_07089_),
    .B1(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__nor2_1 _14563_ (.A(_07297_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__and2b_1 _14564_ (.A_N(_07295_),
    .B(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__and2_1 _14565_ (.A(_07294_),
    .B(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__nor2_1 _14566_ (.A(_07294_),
    .B(_07301_),
    .Y(_07303_));
 sky130_fd_sc_hd__nor2_1 _14567_ (.A(_07302_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__xor2_1 _14568_ (.A(_07297_),
    .B(_07299_),
    .X(_07305_));
 sky130_fd_sc_hd__nand2_1 _14569_ (.A(_07305_),
    .B(_07093_),
    .Y(_07306_));
 sky130_fd_sc_hd__xor2_1 _14570_ (.A(_07295_),
    .B(_07300_),
    .X(_07307_));
 sky130_fd_sc_hd__nand2_1 _14571_ (.A(_07306_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__nand2_1 _14572_ (.A(_07095_),
    .B(_07096_),
    .Y(_07309_));
 sky130_fd_sc_hd__xnor2_1 _14573_ (.A(_07305_),
    .B(_07093_),
    .Y(_07310_));
 sky130_fd_sc_hd__nand2_1 _14574_ (.A(_07309_),
    .B(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__and3_1 _14575_ (.A(_07305_),
    .B(_07095_),
    .C(_07096_),
    .X(_07312_));
 sky130_fd_sc_hd__a221o_1 _14576_ (.A1(_07095_),
    .A2(_07035_),
    .B1(_07043_),
    .B2(_07098_),
    .C1(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__nor2_1 _14577_ (.A(_07295_),
    .B(_07306_),
    .Y(_07314_));
 sky130_fd_sc_hd__a21o_1 _14578_ (.A1(_07311_),
    .A2(_07313_),
    .B1(_07314_),
    .X(_07315_));
 sky130_fd_sc_hd__nand2_1 _14579_ (.A(_07285_),
    .B(_07293_),
    .Y(_07316_));
 sky130_fd_sc_hd__xor2_2 _14580_ (.A(_07273_),
    .B(_07278_),
    .X(_07317_));
 sky130_fd_sc_hd__nand2_1 _14581_ (.A(_07316_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__nand2_1 _14582_ (.A(_07294_),
    .B(_07301_),
    .Y(_07319_));
 sky130_fd_sc_hd__a21oi_1 _14583_ (.A1(_07316_),
    .A2(_07319_),
    .B1(_07317_),
    .Y(_07320_));
 sky130_fd_sc_hd__a41o_1 _14584_ (.A1(_07304_),
    .A2(_07308_),
    .A3(_07315_),
    .A4(_07318_),
    .B1(_07320_),
    .X(_07321_));
 sky130_fd_sc_hd__o21bai_1 _14585_ (.A1(_07279_),
    .A2(_07282_),
    .B1_N(_07281_),
    .Y(_07322_));
 sky130_fd_sc_hd__a21o_1 _14586_ (.A1(_07284_),
    .A2(_07321_),
    .B1(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__and2_1 _14587_ (.A(_06696_),
    .B(_07072_),
    .X(_07324_));
 sky130_fd_sc_hd__or2_1 _14588_ (.A(_07116_),
    .B(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__a21oi_1 _14589_ (.A1(_07131_),
    .A2(_07325_),
    .B1(_07206_),
    .Y(_07326_));
 sky130_fd_sc_hd__a21oi_1 _14590_ (.A1(_07203_),
    .A2(_07210_),
    .B1(_07154_),
    .Y(_07327_));
 sky130_fd_sc_hd__xnor2_1 _14591_ (.A(_07326_),
    .B(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__nor2_1 _14592_ (.A(_07213_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand2_1 _14593_ (.A(_07213_),
    .B(_07328_),
    .Y(_07330_));
 sky130_fd_sc_hd__and2b_1 _14594_ (.A_N(_07329_),
    .B(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__and2_1 _14595_ (.A(_07216_),
    .B(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__nor2_1 _14596_ (.A(_07216_),
    .B(_07331_),
    .Y(_07333_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(_07332_),
    .B(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__a31o_1 _14598_ (.A1(_07218_),
    .A2(_07323_),
    .A3(_07334_),
    .B1(_07332_),
    .X(_07335_));
 sky130_fd_sc_hd__a211o_1 _14599_ (.A1(_07218_),
    .A2(_07323_),
    .B1(_07331_),
    .C1(_07216_),
    .X(_07336_));
 sky130_fd_sc_hd__or3b_1 _14600_ (.A(_07107_),
    .B(_07335_),
    .C_N(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__and2b_1 _14601_ (.A_N(_07327_),
    .B(_07326_),
    .X(_07338_));
 sky130_fd_sc_hd__a2bb2o_1 _14602_ (.A1_N(_07149_),
    .A2_N(_07324_),
    .B1(_06176_),
    .B2(_07116_),
    .X(_07339_));
 sky130_fd_sc_hd__o21ai_1 _14603_ (.A1(_07206_),
    .A2(_07338_),
    .B1(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__or3_1 _14604_ (.A(_07206_),
    .B(_07339_),
    .C(_07338_),
    .X(_07341_));
 sky130_fd_sc_hd__and2_1 _14605_ (.A(_07340_),
    .B(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__nand3b_1 _14606_ (.A_N(_07329_),
    .B(_07330_),
    .C(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__a21oi_1 _14607_ (.A1(_07218_),
    .A2(_07323_),
    .B1(_07216_),
    .Y(_07344_));
 sky130_fd_sc_hd__xnor2_1 _14608_ (.A(_07330_),
    .B(_07342_),
    .Y(_07345_));
 sky130_fd_sc_hd__a311o_1 _14609_ (.A1(_07218_),
    .A2(_07323_),
    .A3(_07334_),
    .B1(_07332_),
    .C1(_07345_),
    .X(_07346_));
 sky130_fd_sc_hd__o211ai_2 _14610_ (.A1(_07343_),
    .A2(_07344_),
    .B1(_07346_),
    .C1(_07107_),
    .Y(_07347_));
 sky130_fd_sc_hd__nand3_1 _14611_ (.A(_07106_),
    .B(_07337_),
    .C(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__xor2_1 _14612_ (.A(_07218_),
    .B(_07323_),
    .X(_07349_));
 sky130_fd_sc_hd__xor2_1 _14613_ (.A(_07284_),
    .B(_07321_),
    .X(_07350_));
 sky130_fd_sc_hd__and2_1 _14614_ (.A(_05793_),
    .B(_07350_),
    .X(_07351_));
 sky130_fd_sc_hd__a21o_1 _14615_ (.A1(_07107_),
    .A2(_07349_),
    .B1(_07351_),
    .X(_07352_));
 sky130_fd_sc_hd__or2_1 _14616_ (.A(_05931_),
    .B(_07352_),
    .X(_07353_));
 sky130_fd_sc_hd__and3_1 _14617_ (.A(_07304_),
    .B(_07308_),
    .C(_07315_),
    .X(_07354_));
 sky130_fd_sc_hd__a21oi_1 _14618_ (.A1(_07308_),
    .A2(_07315_),
    .B1(_07304_),
    .Y(_07355_));
 sky130_fd_sc_hd__nor2_1 _14619_ (.A(_07354_),
    .B(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__and2_1 _14620_ (.A(_05793_),
    .B(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__xnor2_1 _14621_ (.A(_07316_),
    .B(_07317_),
    .Y(_07358_));
 sky130_fd_sc_hd__a31o_1 _14622_ (.A1(_07304_),
    .A2(_07308_),
    .A3(_07315_),
    .B1(_07302_),
    .X(_07359_));
 sky130_fd_sc_hd__xnor2_1 _14623_ (.A(_07358_),
    .B(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__and2_1 _14624_ (.A(_05893_),
    .B(_07360_),
    .X(_07361_));
 sky130_fd_sc_hd__or2_1 _14625_ (.A(_07357_),
    .B(_07361_),
    .X(_07362_));
 sky130_fd_sc_hd__a21oi_1 _14626_ (.A1(_07095_),
    .A2(_07035_),
    .B1(_07099_),
    .Y(_07363_));
 sky130_fd_sc_hd__a21oi_1 _14627_ (.A1(_07309_),
    .A2(_07310_),
    .B1(_07312_),
    .Y(_07364_));
 sky130_fd_sc_hd__xnor2_1 _14628_ (.A(_07363_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__nand2_1 _14629_ (.A(_05793_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__and2_1 _14630_ (.A(_07306_),
    .B(_07307_),
    .X(_07367_));
 sky130_fd_sc_hd__o211ai_1 _14631_ (.A1(_07314_),
    .A2(_07367_),
    .B1(_07311_),
    .C1(_07313_),
    .Y(_07368_));
 sky130_fd_sc_hd__o21ai_1 _14632_ (.A1(_07367_),
    .A2(_07315_),
    .B1(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__nand2_1 _14633_ (.A(_05893_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_1 _14634_ (.A(_07366_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__or2_1 _14635_ (.A(_05931_),
    .B(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__o211a_1 _14636_ (.A1(_05779_),
    .A2(_07362_),
    .B1(_07372_),
    .C1(_05892_),
    .X(_07373_));
 sky130_fd_sc_hd__a31o_1 _14637_ (.A1(_05741_),
    .A2(_07348_),
    .A3(_07353_),
    .B1(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__buf_2 _14638_ (.A(_05932_),
    .X(_07375_));
 sky130_fd_sc_hd__a32o_1 _14639_ (.A1(_05742_),
    .A2(_05755_),
    .A3(_07105_),
    .B1(_07374_),
    .B2(_07375_),
    .X(_07376_));
 sky130_fd_sc_hd__and3_1 _14640_ (.A(_07106_),
    .B(_07107_),
    .C(_07041_),
    .X(_07377_));
 sky130_fd_sc_hd__buf_2 _14641_ (.A(_05793_),
    .X(_07378_));
 sky130_fd_sc_hd__nand2_1 _14642_ (.A(_07378_),
    .B(_07349_),
    .Y(_07379_));
 sky130_fd_sc_hd__or3b_1 _14643_ (.A(_07378_),
    .B(_07335_),
    .C_N(_07336_),
    .X(_07380_));
 sky130_fd_sc_hd__mux2_1 _14644_ (.A0(_07350_),
    .A1(_07360_),
    .S(_05793_),
    .X(_07381_));
 sky130_fd_sc_hd__nor2_1 _14645_ (.A(_05931_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__a31o_1 _14646_ (.A1(_07106_),
    .A2(_07379_),
    .A3(_07380_),
    .B1(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__nor2_1 _14647_ (.A(_05893_),
    .B(_07101_),
    .Y(_07384_));
 sky130_fd_sc_hd__and2_1 _14648_ (.A(_05893_),
    .B(_07365_),
    .X(_07385_));
 sky130_fd_sc_hd__or2_1 _14649_ (.A(_07384_),
    .B(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__nand2_1 _14650_ (.A(_05793_),
    .B(_07369_),
    .Y(_07387_));
 sky130_fd_sc_hd__a21bo_1 _14651_ (.A1(_07107_),
    .A2(_07356_),
    .B1_N(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(_07386_),
    .A1(_07388_),
    .S(_05931_),
    .X(_07389_));
 sky130_fd_sc_hd__nor2_1 _14653_ (.A(_05741_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__a21oi_1 _14654_ (.A1(_05741_),
    .A2(_07383_),
    .B1(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__a32o_1 _14655_ (.A1(_05742_),
    .A2(_05755_),
    .A3(_07377_),
    .B1(_07391_),
    .B2(_07375_),
    .X(_07392_));
 sky130_fd_sc_hd__or2_1 _14656_ (.A(_05703_),
    .B(_05928_),
    .X(_07393_));
 sky130_fd_sc_hd__buf_2 _14657_ (.A(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(_07352_),
    .A1(_07362_),
    .S(_05779_),
    .X(_07395_));
 sky130_fd_sc_hd__clkinv_2 _14659_ (.A(_07103_),
    .Y(_07396_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(_07371_),
    .A1(_07396_),
    .S(_05779_),
    .X(_07397_));
 sky130_fd_sc_hd__or2_1 _14661_ (.A(_05741_),
    .B(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__o211a_1 _14662_ (.A1(_05892_),
    .A2(_07395_),
    .B1(_07398_),
    .C1(_07375_),
    .X(_07399_));
 sky130_fd_sc_hd__mux2_1 _14663_ (.A0(_07388_),
    .A1(_07381_),
    .S(_05931_),
    .X(_07400_));
 sky130_fd_sc_hd__and2_1 _14664_ (.A(_05893_),
    .B(_07041_),
    .X(_07401_));
 sky130_fd_sc_hd__mux2_1 _14665_ (.A0(_07386_),
    .A1(_07401_),
    .S(_05779_),
    .X(_07402_));
 sky130_fd_sc_hd__mux2_1 _14666_ (.A0(_07400_),
    .A1(_07402_),
    .S(_05892_),
    .X(_07403_));
 sky130_fd_sc_hd__nand2_1 _14667_ (.A(_07375_),
    .B(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__or3b_1 _14668_ (.A(_07394_),
    .B(_07399_),
    .C_N(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__or3_1 _14669_ (.A(_07376_),
    .B(_07392_),
    .C(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__and4_1 _14670_ (.A(_07218_),
    .B(_07323_),
    .C(_07345_),
    .D(_07334_),
    .X(_07407_));
 sky130_fd_sc_hd__a21o_1 _14671_ (.A1(_07213_),
    .A2(_07328_),
    .B1(_07332_),
    .X(_07408_));
 sky130_fd_sc_hd__nand2_1 _14672_ (.A(_07342_),
    .B(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__inv_2 _14673_ (.A(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__nor2_1 _14674_ (.A(_06239_),
    .B(_07149_),
    .Y(_07411_));
 sky130_fd_sc_hd__o211a_1 _14675_ (.A1(_06724_),
    .A2(_06761_),
    .B1(_07411_),
    .C1(_07340_),
    .X(_07412_));
 sky130_fd_sc_hd__o21ba_2 _14676_ (.A1(_07407_),
    .A2(_07410_),
    .B1_N(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__and3b_1 _14677_ (.A_N(_07407_),
    .B(_07409_),
    .C(_07412_),
    .X(_07414_));
 sky130_fd_sc_hd__nor3_1 _14678_ (.A(_07378_),
    .B(_07413_),
    .C(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__o211a_1 _14679_ (.A1(_07343_),
    .A2(_07344_),
    .B1(_07346_),
    .C1(_07378_),
    .X(_07416_));
 sky130_fd_sc_hd__a211o_1 _14680_ (.A1(_07378_),
    .A2(_07413_),
    .B1(_06239_),
    .C1(_05779_),
    .X(_07417_));
 sky130_fd_sc_hd__o311a_1 _14681_ (.A1(_07106_),
    .A2(_07415_),
    .A3(_07416_),
    .B1(_07417_),
    .C1(_05892_),
    .X(_07418_));
 sky130_fd_sc_hd__nand2_2 _14682_ (.A(_07107_),
    .B(_07413_),
    .Y(_07419_));
 sky130_fd_sc_hd__or3_2 _14683_ (.A(_07107_),
    .B(_07413_),
    .C(_07414_),
    .X(_07420_));
 sky130_fd_sc_hd__a211o_1 _14684_ (.A1(_07419_),
    .A2(_07420_),
    .B1(_05741_),
    .C1(_07106_),
    .X(_07421_));
 sky130_fd_sc_hd__nand2_1 _14685_ (.A(_07394_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__and3_1 _14686_ (.A(_05779_),
    .B(_07337_),
    .C(_07347_),
    .X(_07423_));
 sky130_fd_sc_hd__a311oi_2 _14687_ (.A1(_07106_),
    .A2(_07419_),
    .A3(_07420_),
    .B1(_07423_),
    .C1(_05742_),
    .Y(_07424_));
 sky130_fd_sc_hd__a21oi_1 _14688_ (.A1(_07378_),
    .A2(_07413_),
    .B1(_06239_),
    .Y(_07425_));
 sky130_fd_sc_hd__or2_1 _14689_ (.A(_07106_),
    .B(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__o211ai_1 _14690_ (.A1(_07343_),
    .A2(_07344_),
    .B1(_07346_),
    .C1(_07378_),
    .Y(_07427_));
 sky130_fd_sc_hd__o31a_1 _14691_ (.A1(_07378_),
    .A2(_07413_),
    .A3(_07414_),
    .B1(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__a21o_1 _14692_ (.A1(_07379_),
    .A2(_07380_),
    .B1(_05931_),
    .X(_07429_));
 sky130_fd_sc_hd__o211a_1 _14693_ (.A1(_05779_),
    .A2(_07428_),
    .B1(_07429_),
    .C1(_05892_),
    .X(_07430_));
 sky130_fd_sc_hd__a21o_1 _14694_ (.A1(_05742_),
    .A2(_07426_),
    .B1(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__or4b_1 _14695_ (.A(_07418_),
    .B(_07422_),
    .C(_07424_),
    .D_N(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__clkbuf_4 _14696_ (.A(_07375_),
    .X(_07433_));
 sky130_fd_sc_hd__nand2_1 _14697_ (.A(_07394_),
    .B(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__a311o_1 _14698_ (.A1(_07106_),
    .A2(_07419_),
    .A3(_07420_),
    .B1(_07423_),
    .C1(_05892_),
    .X(_07435_));
 sky130_fd_sc_hd__nand2_1 _14699_ (.A(_05892_),
    .B(_07395_),
    .Y(_07436_));
 sky130_fd_sc_hd__nand2_1 _14700_ (.A(_05741_),
    .B(_07397_),
    .Y(_07437_));
 sky130_fd_sc_hd__and2_1 _14701_ (.A(_05963_),
    .B(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__a31o_1 _14702_ (.A1(_07375_),
    .A2(_07435_),
    .A3(_07436_),
    .B1(_07438_),
    .X(_07439_));
 sky130_fd_sc_hd__o311ai_2 _14703_ (.A1(_07106_),
    .A2(_07415_),
    .A3(_07416_),
    .B1(_07417_),
    .C1(_05742_),
    .Y(_07440_));
 sky130_fd_sc_hd__or2_1 _14704_ (.A(_05741_),
    .B(_07383_),
    .X(_07441_));
 sky130_fd_sc_hd__a22o_1 _14705_ (.A1(_05894_),
    .A2(_07041_),
    .B1(_07389_),
    .B2(_05741_),
    .X(_07442_));
 sky130_fd_sc_hd__nor2_1 _14706_ (.A(_07375_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__a31o_1 _14707_ (.A1(_07375_),
    .A2(_07440_),
    .A3(_07441_),
    .B1(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__o211a_1 _14708_ (.A1(_05779_),
    .A2(_07428_),
    .B1(_07429_),
    .C1(_05742_),
    .X(_07445_));
 sky130_fd_sc_hd__nor2_1 _14709_ (.A(_05742_),
    .B(_07400_),
    .Y(_07446_));
 sky130_fd_sc_hd__nand2_1 _14710_ (.A(_05741_),
    .B(_07402_),
    .Y(_07447_));
 sky130_fd_sc_hd__or2_1 _14711_ (.A(_07375_),
    .B(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__o31a_1 _14712_ (.A1(_05963_),
    .A2(_07445_),
    .A3(_07446_),
    .B1(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__o21ai_1 _14713_ (.A1(_05779_),
    .A2(_07362_),
    .B1(_07372_),
    .Y(_07450_));
 sky130_fd_sc_hd__nand2_1 _14714_ (.A(_07348_),
    .B(_07353_),
    .Y(_07451_));
 sky130_fd_sc_hd__a21o_1 _14715_ (.A1(_07419_),
    .A2(_07420_),
    .B1(_07106_),
    .X(_07452_));
 sky130_fd_sc_hd__mux4_2 _14716_ (.A0(_07104_),
    .A1(_07450_),
    .A2(_07451_),
    .A3(_07452_),
    .S0(_05742_),
    .S1(_07375_),
    .X(_07453_));
 sky130_fd_sc_hd__nand4_1 _14717_ (.A(_07439_),
    .B(_07444_),
    .C(_07449_),
    .D(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__a32o_4 _14718_ (.A1(_07406_),
    .A2(_07432_),
    .A3(_07434_),
    .B1(_07454_),
    .B2(_05929_),
    .X(_07455_));
 sky130_fd_sc_hd__buf_4 _14719_ (.A(_07455_),
    .X(_07456_));
 sky130_fd_sc_hd__inv_2 _14720_ (.A(_07431_),
    .Y(_07457_));
 sky130_fd_sc_hd__mux2_1 _14721_ (.A0(_07403_),
    .A1(_07457_),
    .S(_07433_),
    .X(_07458_));
 sky130_fd_sc_hd__buf_4 _14722_ (.A(_05871_),
    .X(_07459_));
 sky130_fd_sc_hd__mux2_1 _14723_ (.A0(_07456_),
    .A1(_07458_),
    .S(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__clkbuf_4 _14724_ (.A(_05188_),
    .X(_07461_));
 sky130_fd_sc_hd__mux2_1 _14725_ (.A0(\rbzero.wall_tracer.stepDistY[-12] ),
    .A1(_07460_),
    .S(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__clkbuf_1 _14726_ (.A(_07462_),
    .X(_00419_));
 sky130_fd_sc_hd__o21a_1 _14727_ (.A1(_05892_),
    .A2(_07395_),
    .B1(_07398_),
    .X(_07463_));
 sky130_fd_sc_hd__mux2_1 _14728_ (.A0(_07463_),
    .A1(_07424_),
    .S(_07433_),
    .X(_07464_));
 sky130_fd_sc_hd__mux2_2 _14729_ (.A0(_07456_),
    .A1(_07464_),
    .S(_07459_),
    .X(_07465_));
 sky130_fd_sc_hd__mux2_1 _14730_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_07465_),
    .S(_07461_),
    .X(_07466_));
 sky130_fd_sc_hd__clkbuf_1 _14731_ (.A(_07466_),
    .X(_00420_));
 sky130_fd_sc_hd__and2_1 _14732_ (.A(_05834_),
    .B(_07455_),
    .X(_07467_));
 sky130_fd_sc_hd__clkbuf_4 _14733_ (.A(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__a21o_1 _14734_ (.A1(_07378_),
    .A2(_07413_),
    .B1(_07415_),
    .X(_07469_));
 sky130_fd_sc_hd__nand2_1 _14735_ (.A(_07380_),
    .B(_07427_),
    .Y(_07470_));
 sky130_fd_sc_hd__mux2_1 _14736_ (.A0(_07469_),
    .A1(_07470_),
    .S(_05952_),
    .X(_07471_));
 sky130_fd_sc_hd__a21o_1 _14737_ (.A1(_05844_),
    .A2(_07471_),
    .B1(_06239_),
    .X(_07472_));
 sky130_fd_sc_hd__buf_2 _14738_ (.A(_05844_),
    .X(_07473_));
 sky130_fd_sc_hd__and2_1 _14739_ (.A(_07378_),
    .B(_07360_),
    .X(_07474_));
 sky130_fd_sc_hd__a21oi_1 _14740_ (.A1(_07107_),
    .A2(_07356_),
    .B1(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__a21boi_1 _14741_ (.A1(_07107_),
    .A2(_07350_),
    .B1_N(_07379_),
    .Y(_07476_));
 sky130_fd_sc_hd__clkbuf_4 _14742_ (.A(_05807_),
    .X(_07477_));
 sky130_fd_sc_hd__mux2_1 _14743_ (.A0(_07475_),
    .A1(_07476_),
    .S(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__or2b_1 _14744_ (.A(_07385_),
    .B_N(_07387_),
    .X(_07479_));
 sky130_fd_sc_hd__o211a_1 _14745_ (.A1(_07384_),
    .A2(_07401_),
    .B1(_05844_),
    .C1(_05952_),
    .X(_07480_));
 sky130_fd_sc_hd__a311o_1 _14746_ (.A1(_05844_),
    .A2(_07477_),
    .A3(_07479_),
    .B1(_07480_),
    .C1(_05800_),
    .X(_07481_));
 sky130_fd_sc_hd__o21bai_1 _14747_ (.A1(_07473_),
    .A2(_07478_),
    .B1_N(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__o211a_1 _14748_ (.A1(_05814_),
    .A2(_07472_),
    .B1(_07482_),
    .C1(_07459_),
    .X(_07483_));
 sky130_fd_sc_hd__or2_1 _14749_ (.A(_07468_),
    .B(_07483_),
    .X(_07484_));
 sky130_fd_sc_hd__mux2_1 _14750_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_07484_),
    .S(_07461_),
    .X(_07485_));
 sky130_fd_sc_hd__clkbuf_1 _14751_ (.A(_07485_),
    .X(_00421_));
 sky130_fd_sc_hd__buf_4 _14752_ (.A(_05834_),
    .X(_07486_));
 sky130_fd_sc_hd__buf_4 _14753_ (.A(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__nor2_1 _14754_ (.A(_05794_),
    .B(_07104_),
    .Y(_07488_));
 sky130_fd_sc_hd__a21bo_1 _14755_ (.A1(_07107_),
    .A2(_07349_),
    .B1_N(_07337_),
    .X(_07489_));
 sky130_fd_sc_hd__nor2_1 _14756_ (.A(_07351_),
    .B(_07361_),
    .Y(_07490_));
 sky130_fd_sc_hd__nor2_1 _14757_ (.A(_07477_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__a21oi_1 _14758_ (.A1(_07477_),
    .A2(_07489_),
    .B1(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__and2b_1 _14759_ (.A_N(_07357_),
    .B(_07370_),
    .X(_07493_));
 sky130_fd_sc_hd__and4b_1 _14760_ (.A_N(_07102_),
    .B(_05952_),
    .C(_05844_),
    .D(_07366_),
    .X(_07494_));
 sky130_fd_sc_hd__a31o_1 _14761_ (.A1(_07473_),
    .A2(_07477_),
    .A3(_07493_),
    .B1(_07494_),
    .X(_07495_));
 sky130_fd_sc_hd__a21o_1 _14762_ (.A1(_05884_),
    .A2(_07492_),
    .B1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__clkinv_2 _14763_ (.A(_07419_),
    .Y(_07497_));
 sky130_fd_sc_hd__nand2_1 _14764_ (.A(_07420_),
    .B(_07347_),
    .Y(_07498_));
 sky130_fd_sc_hd__mux2_1 _14765_ (.A0(_07497_),
    .A1(_07498_),
    .S(_05952_),
    .X(_07499_));
 sky130_fd_sc_hd__a21oi_1 _14766_ (.A1(_07473_),
    .A2(_07499_),
    .B1(_05814_),
    .Y(_07500_));
 sky130_fd_sc_hd__a211oi_1 _14767_ (.A1(_05814_),
    .A2(_07496_),
    .B1(_07500_),
    .C1(_07486_),
    .Y(_07501_));
 sky130_fd_sc_hd__a211o_1 _14768_ (.A1(_07487_),
    .A2(_07455_),
    .B1(_07488_),
    .C1(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__mux2_1 _14769_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_07502_),
    .S(_07461_),
    .X(_07503_));
 sky130_fd_sc_hd__clkbuf_1 _14770_ (.A(_07503_),
    .X(_00422_));
 sky130_fd_sc_hd__and3_1 _14771_ (.A(_05844_),
    .B(_05952_),
    .C(_07469_),
    .X(_07504_));
 sky130_fd_sc_hd__or2_1 _14772_ (.A(_05814_),
    .B(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__nor2_1 _14773_ (.A(_07477_),
    .B(_07476_),
    .Y(_07506_));
 sky130_fd_sc_hd__a21oi_1 _14774_ (.A1(_07477_),
    .A2(_07470_),
    .B1(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__nor2_1 _14775_ (.A(_07477_),
    .B(_07479_),
    .Y(_07508_));
 sky130_fd_sc_hd__a211o_1 _14776_ (.A1(_07477_),
    .A2(_07475_),
    .B1(_07508_),
    .C1(_05884_),
    .X(_07509_));
 sky130_fd_sc_hd__o211ai_1 _14777_ (.A1(_07473_),
    .A2(_07507_),
    .B1(_07509_),
    .C1(_05814_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand2_1 _14778_ (.A(_07486_),
    .B(_07433_),
    .Y(_07511_));
 sky130_fd_sc_hd__nor2_1 _14779_ (.A(_07511_),
    .B(_07447_),
    .Y(_07512_));
 sky130_fd_sc_hd__a31o_1 _14780_ (.A1(_07459_),
    .A2(_07505_),
    .A3(_07510_),
    .B1(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__a21oi_4 _14781_ (.A1(_07487_),
    .A2(_07456_),
    .B1(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__nor2_1 _14782_ (.A(\rbzero.wall_tracer.stepDistY[-8] ),
    .B(_00004_),
    .Y(_07515_));
 sky130_fd_sc_hd__a21oi_1 _14783_ (.A1(_00004_),
    .A2(_07514_),
    .B1(_07515_),
    .Y(_00423_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(_07498_),
    .A1(_07489_),
    .S(_05952_),
    .X(_07516_));
 sky130_fd_sc_hd__mux2_1 _14785_ (.A0(_07490_),
    .A1(_07493_),
    .S(_05952_),
    .X(_07517_));
 sky130_fd_sc_hd__nor2_1 _14786_ (.A(_05884_),
    .B(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__a211o_1 _14787_ (.A1(_05884_),
    .A2(_07516_),
    .B1(_07518_),
    .C1(_05800_),
    .X(_07519_));
 sky130_fd_sc_hd__or3_1 _14788_ (.A(_05884_),
    .B(_07477_),
    .C(_07419_),
    .X(_07520_));
 sky130_fd_sc_hd__nand2_1 _14789_ (.A(_05800_),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__and3_1 _14790_ (.A(_07459_),
    .B(_07519_),
    .C(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__nor2_1 _14791_ (.A(_07511_),
    .B(_07437_),
    .Y(_07523_));
 sky130_fd_sc_hd__a211oi_4 _14792_ (.A1(_07487_),
    .A2(_07456_),
    .B1(_07522_),
    .C1(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__nor2_1 _14793_ (.A(\rbzero.wall_tracer.stepDistY[-7] ),
    .B(_00004_),
    .Y(_07525_));
 sky130_fd_sc_hd__a21oi_1 _14794_ (.A1(_00004_),
    .A2(_07524_),
    .B1(_07525_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _14795_ (.A(_07473_),
    .B(_07478_),
    .Y(_07526_));
 sky130_fd_sc_hd__nor2_2 _14796_ (.A(_05834_),
    .B(_05800_),
    .Y(_07527_));
 sky130_fd_sc_hd__o211a_1 _14797_ (.A1(_07473_),
    .A2(_07471_),
    .B1(_07526_),
    .C1(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__a31o_1 _14798_ (.A1(_07486_),
    .A2(_07433_),
    .A3(_07442_),
    .B1(_07528_),
    .X(_07529_));
 sky130_fd_sc_hd__a21oi_4 _14799_ (.A1(_07487_),
    .A2(_07456_),
    .B1(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__nor2_1 _14800_ (.A(\rbzero.wall_tracer.stepDistY[-6] ),
    .B(_07461_),
    .Y(_07531_));
 sky130_fd_sc_hd__a21oi_1 _14801_ (.A1(_00004_),
    .A2(_07530_),
    .B1(_07531_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _14802_ (.A(_07473_),
    .B(_07492_),
    .Y(_07532_));
 sky130_fd_sc_hd__o211a_1 _14803_ (.A1(_07473_),
    .A2(_07499_),
    .B1(_07532_),
    .C1(_07527_),
    .X(_07533_));
 sky130_fd_sc_hd__mux2_1 _14804_ (.A0(_07104_),
    .A1(_07450_),
    .S(_05742_),
    .X(_07534_));
 sky130_fd_sc_hd__nor2_1 _14805_ (.A(_07511_),
    .B(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__a211oi_4 _14806_ (.A1(_07487_),
    .A2(_07456_),
    .B1(_07533_),
    .C1(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__nor2_1 _14807_ (.A(\rbzero.wall_tracer.stepDistY[-5] ),
    .B(_07461_),
    .Y(_07537_));
 sky130_fd_sc_hd__a21oi_1 _14808_ (.A1(_00004_),
    .A2(_07536_),
    .B1(_07537_),
    .Y(_00426_));
 sky130_fd_sc_hd__nor2_1 _14809_ (.A(_05884_),
    .B(_07507_),
    .Y(_07538_));
 sky130_fd_sc_hd__a31o_1 _14810_ (.A1(_05884_),
    .A2(_05952_),
    .A3(_07469_),
    .B1(_07538_),
    .X(_07539_));
 sky130_fd_sc_hd__nor2_1 _14811_ (.A(_07459_),
    .B(_07404_),
    .Y(_07540_));
 sky130_fd_sc_hd__a221o_4 _14812_ (.A1(_07486_),
    .A2(_07455_),
    .B1(_07539_),
    .B2(_07527_),
    .C1(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__mux2_1 _14813_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_07541_),
    .S(_07461_),
    .X(_07542_));
 sky130_fd_sc_hd__clkbuf_1 _14814_ (.A(_07542_),
    .X(_00427_));
 sky130_fd_sc_hd__a22o_1 _14815_ (.A1(_05894_),
    .A2(_07413_),
    .B1(_07516_),
    .B2(_07473_),
    .X(_07543_));
 sky130_fd_sc_hd__a22o_1 _14816_ (.A1(_07486_),
    .A2(_07399_),
    .B1(_07543_),
    .B2(_07527_),
    .X(_07544_));
 sky130_fd_sc_hd__a21o_1 _14817_ (.A1(_07487_),
    .A2(_07456_),
    .B1(_07544_),
    .X(_07545_));
 sky130_fd_sc_hd__buf_4 _14818_ (.A(_05188_),
    .X(_07546_));
 sky130_fd_sc_hd__mux2_1 _14819_ (.A0(\rbzero.wall_tracer.stepDistY[-3] ),
    .A1(_07545_),
    .S(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__clkbuf_1 _14820_ (.A(_07547_),
    .X(_00428_));
 sky130_fd_sc_hd__a22o_1 _14821_ (.A1(_05834_),
    .A2(_07392_),
    .B1(_07472_),
    .B2(_07527_),
    .X(_07548_));
 sky130_fd_sc_hd__a21oi_4 _14822_ (.A1(_07486_),
    .A2(_07455_),
    .B1(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(\rbzero.wall_tracer.stepDistY[-2] ),
    .B(_07461_),
    .Y(_07550_));
 sky130_fd_sc_hd__a21oi_1 _14824_ (.A1(_00004_),
    .A2(_07549_),
    .B1(_07550_),
    .Y(_00429_));
 sky130_fd_sc_hd__a32o_2 _14825_ (.A1(_07473_),
    .A2(_07527_),
    .A3(_07499_),
    .B1(_07376_),
    .B2(_05834_),
    .X(_07551_));
 sky130_fd_sc_hd__a21oi_4 _14826_ (.A1(_07486_),
    .A2(_07455_),
    .B1(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__nor2_1 _14827_ (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .B(_07461_),
    .Y(_07553_));
 sky130_fd_sc_hd__a21oi_1 _14828_ (.A1(_00004_),
    .A2(_07552_),
    .B1(_07553_),
    .Y(_00430_));
 sky130_fd_sc_hd__o2bb2a_1 _14829_ (.A1_N(_07527_),
    .A2_N(_07504_),
    .B1(_07449_),
    .B2(_07459_),
    .X(_07554_));
 sky130_fd_sc_hd__a21boi_4 _14830_ (.A1(_07486_),
    .A2(_07455_),
    .B1_N(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__nor2_1 _14831_ (.A(\rbzero.wall_tracer.stepDistY[0] ),
    .B(_07461_),
    .Y(_07556_));
 sky130_fd_sc_hd__a21oi_1 _14832_ (.A1(_00004_),
    .A2(_07555_),
    .B1(_07556_),
    .Y(_00431_));
 sky130_fd_sc_hd__nor2_1 _14833_ (.A(_07459_),
    .B(_07439_),
    .Y(_07557_));
 sky130_fd_sc_hd__or3_1 _14834_ (.A(_05834_),
    .B(_05800_),
    .C(_07520_),
    .X(_07558_));
 sky130_fd_sc_hd__or3b_1 _14835_ (.A(_07468_),
    .B(_07557_),
    .C_N(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__clkbuf_4 _14836_ (.A(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__mux2_1 _14837_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_07560_),
    .S(_07546_),
    .X(_07561_));
 sky130_fd_sc_hd__clkbuf_1 _14838_ (.A(_07561_),
    .X(_00432_));
 sky130_fd_sc_hd__o21bai_4 _14839_ (.A1(_07459_),
    .A2(_07444_),
    .B1_N(_07468_),
    .Y(_07562_));
 sky130_fd_sc_hd__mux2_1 _14840_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_07562_),
    .S(_07546_),
    .X(_07563_));
 sky130_fd_sc_hd__clkbuf_1 _14841_ (.A(_07563_),
    .X(_00433_));
 sky130_fd_sc_hd__o21bai_4 _14842_ (.A1(_07459_),
    .A2(_07453_),
    .B1_N(_07468_),
    .Y(_07564_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_07564_),
    .S(_07546_),
    .X(_07565_));
 sky130_fd_sc_hd__clkbuf_1 _14844_ (.A(_07565_),
    .X(_00434_));
 sky130_fd_sc_hd__o31a_2 _14845_ (.A1(_05929_),
    .A2(_07456_),
    .A3(_07458_),
    .B1(_07487_),
    .X(_07566_));
 sky130_fd_sc_hd__mux2_1 _14846_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_07566_),
    .S(_07546_),
    .X(_07567_));
 sky130_fd_sc_hd__clkbuf_1 _14847_ (.A(_07567_),
    .X(_00435_));
 sky130_fd_sc_hd__a21o_2 _14848_ (.A1(_07394_),
    .A2(_07464_),
    .B1(_07468_),
    .X(_07568_));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_07568_),
    .S(_07546_),
    .X(_07569_));
 sky130_fd_sc_hd__clkbuf_1 _14850_ (.A(_07569_),
    .X(_00436_));
 sky130_fd_sc_hd__a2111oi_1 _14851_ (.A1(_05742_),
    .A2(_07383_),
    .B1(_07390_),
    .C1(_05736_),
    .D1(_05737_),
    .Y(_07570_));
 sky130_fd_sc_hd__a311o_4 _14852_ (.A1(_07394_),
    .A2(_07433_),
    .A3(_07418_),
    .B1(_07468_),
    .C1(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_07571_),
    .S(_07546_),
    .X(_07572_));
 sky130_fd_sc_hd__clkbuf_1 _14854_ (.A(_07572_),
    .X(_00437_));
 sky130_fd_sc_hd__nand2_1 _14855_ (.A(_07433_),
    .B(_07421_),
    .Y(_07573_));
 sky130_fd_sc_hd__o211ai_4 _14856_ (.A1(_07433_),
    .A2(_07374_),
    .B1(_07573_),
    .C1(_07394_),
    .Y(_07574_));
 sky130_fd_sc_hd__nand2b_4 _14857_ (.A_N(_07468_),
    .B(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__mux2_1 _14858_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_07575_),
    .S(_07546_),
    .X(_07576_));
 sky130_fd_sc_hd__clkbuf_1 _14859_ (.A(_07576_),
    .X(_00438_));
 sky130_fd_sc_hd__nor3_1 _14860_ (.A(_07433_),
    .B(_07445_),
    .C(_07446_),
    .Y(_07577_));
 sky130_fd_sc_hd__o21ai_1 _14861_ (.A1(_05902_),
    .A2(_07426_),
    .B1(_07394_),
    .Y(_07578_));
 sky130_fd_sc_hd__o31a_2 _14862_ (.A1(_07456_),
    .A2(_07577_),
    .A3(_07578_),
    .B1(_07487_),
    .X(_07579_));
 sky130_fd_sc_hd__mux2_1 _14863_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_07579_),
    .S(_07546_),
    .X(_07580_));
 sky130_fd_sc_hd__clkbuf_1 _14864_ (.A(_07580_),
    .X(_00439_));
 sky130_fd_sc_hd__a21oi_1 _14865_ (.A1(_07435_),
    .A2(_07436_),
    .B1(_07433_),
    .Y(_07581_));
 sky130_fd_sc_hd__o31a_2 _14866_ (.A1(_05929_),
    .A2(_07456_),
    .A3(_07581_),
    .B1(_07487_),
    .X(_07582_));
 sky130_fd_sc_hd__mux2_1 _14867_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_07582_),
    .S(_07546_),
    .X(_07583_));
 sky130_fd_sc_hd__clkbuf_1 _14868_ (.A(_07583_),
    .X(_00440_));
 sky130_fd_sc_hd__and3_1 _14869_ (.A(_07394_),
    .B(_07440_),
    .C(_07441_),
    .X(_07584_));
 sky130_fd_sc_hd__or3_2 _14870_ (.A(_05737_),
    .B(_05736_),
    .C(_07584_),
    .X(_07585_));
 sky130_fd_sc_hd__or2b_1 _14871_ (.A(_07468_),
    .B_N(_07585_),
    .X(_07586_));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_07586_),
    .S(_05188_),
    .X(_07587_));
 sky130_fd_sc_hd__clkbuf_1 _14873_ (.A(_07587_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _14874_ (.A0(_07452_),
    .A1(_07451_),
    .S(_05892_),
    .X(_07588_));
 sky130_fd_sc_hd__nor4_4 _14875_ (.A(_05737_),
    .B(_05736_),
    .C(_07588_),
    .D(_07468_),
    .Y(_07589_));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(\rbzero.wall_tracer.stepDistY[11] ),
    .A1(_07589_),
    .S(_05188_),
    .X(_07590_));
 sky130_fd_sc_hd__clkbuf_1 _14877_ (.A(_07590_),
    .X(_00442_));
 sky130_fd_sc_hd__clkbuf_4 _14878_ (.A(_04019_),
    .X(_07591_));
 sky130_fd_sc_hd__buf_4 _14879_ (.A(_05278_),
    .X(_07592_));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(\rbzero.wall_tracer.trackDistY[-12] ),
    .A1(\rbzero.wall_tracer.trackDistX[-12] ),
    .S(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__nor2_2 _14881_ (.A(_03969_),
    .B(_04017_),
    .Y(_07594_));
 sky130_fd_sc_hd__clkbuf_4 _14882_ (.A(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__or2_1 _14883_ (.A(\rbzero.wall_tracer.visualWallDist[-12] ),
    .B(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__o211a_1 _14884_ (.A1(_07591_),
    .A2(_07593_),
    .B1(_07596_),
    .C1(_04039_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _14885_ (.A0(\rbzero.wall_tracer.trackDistY[-11] ),
    .A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .S(_07592_),
    .X(_07597_));
 sky130_fd_sc_hd__inv_2 _14886_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .Y(_07598_));
 sky130_fd_sc_hd__nand2_1 _14887_ (.A(_07598_),
    .B(_04019_),
    .Y(_07599_));
 sky130_fd_sc_hd__o211a_1 _14888_ (.A1(_07591_),
    .A2(_07597_),
    .B1(_07599_),
    .C1(_04039_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _14889_ (.A0(\rbzero.wall_tracer.trackDistY[-10] ),
    .A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .S(_07592_),
    .X(_07600_));
 sky130_fd_sc_hd__buf_4 _14890_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_07601_));
 sky130_fd_sc_hd__clkinv_2 _14891_ (.A(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__nand2_1 _14892_ (.A(_07602_),
    .B(_04019_),
    .Y(_07603_));
 sky130_fd_sc_hd__o211a_1 _14893_ (.A1(_07591_),
    .A2(_07600_),
    .B1(_07603_),
    .C1(_04039_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _14894_ (.A0(\rbzero.wall_tracer.trackDistY[-9] ),
    .A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .S(_07592_),
    .X(_07604_));
 sky130_fd_sc_hd__or2_1 _14895_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_07595_),
    .X(_07605_));
 sky130_fd_sc_hd__o211a_1 _14896_ (.A1(_07591_),
    .A2(_07604_),
    .B1(_07605_),
    .C1(_04039_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _14897_ (.A0(\rbzero.wall_tracer.trackDistY[-8] ),
    .A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .S(_07592_),
    .X(_07606_));
 sky130_fd_sc_hd__or2_1 _14898_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_07595_),
    .X(_07607_));
 sky130_fd_sc_hd__o211a_1 _14899_ (.A1(_07591_),
    .A2(_07606_),
    .B1(_07607_),
    .C1(_04039_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14900_ (.A0(\rbzero.wall_tracer.trackDistY[-7] ),
    .A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .S(_07592_),
    .X(_07608_));
 sky130_fd_sc_hd__or2_1 _14901_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(_07595_),
    .X(_07609_));
 sky130_fd_sc_hd__o211a_1 _14902_ (.A1(_07591_),
    .A2(_07608_),
    .B1(_07609_),
    .C1(_04039_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14903_ (.A0(\rbzero.wall_tracer.trackDistY[-6] ),
    .A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .S(_07592_),
    .X(_07610_));
 sky130_fd_sc_hd__or2_1 _14904_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_07595_),
    .X(_07611_));
 sky130_fd_sc_hd__o211a_1 _14905_ (.A1(_07591_),
    .A2(_07610_),
    .B1(_07611_),
    .C1(_04039_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14906_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .S(_07592_),
    .X(_07612_));
 sky130_fd_sc_hd__or2_1 _14907_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_07595_),
    .X(_07613_));
 sky130_fd_sc_hd__o211a_1 _14908_ (.A1(_07591_),
    .A2(_07612_),
    .B1(_07613_),
    .C1(_04039_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14909_ (.A0(\rbzero.wall_tracer.trackDistY[-4] ),
    .A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .S(_07592_),
    .X(_07614_));
 sky130_fd_sc_hd__or2_1 _14910_ (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .B(_07595_),
    .X(_07615_));
 sky130_fd_sc_hd__o211a_1 _14911_ (.A1(_07591_),
    .A2(_07614_),
    .B1(_07615_),
    .C1(_04039_),
    .X(_00451_));
 sky130_fd_sc_hd__buf_4 _14912_ (.A(_05278_),
    .X(_07616_));
 sky130_fd_sc_hd__mux2_1 _14913_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(\rbzero.wall_tracer.trackDistX[-3] ),
    .S(_07616_),
    .X(_07617_));
 sky130_fd_sc_hd__clkbuf_2 _14914_ (.A(_07594_),
    .X(_07618_));
 sky130_fd_sc_hd__or2_1 _14915_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .B(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__buf_2 _14916_ (.A(_04035_),
    .X(_07620_));
 sky130_fd_sc_hd__o211a_1 _14917_ (.A1(_07591_),
    .A2(_07617_),
    .B1(_07619_),
    .C1(_07620_),
    .X(_00452_));
 sky130_fd_sc_hd__clkbuf_4 _14918_ (.A(_04019_),
    .X(_07621_));
 sky130_fd_sc_hd__mux2_1 _14919_ (.A0(\rbzero.wall_tracer.trackDistY[-2] ),
    .A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .S(_07616_),
    .X(_07622_));
 sky130_fd_sc_hd__or2_1 _14920_ (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .B(_07618_),
    .X(_07623_));
 sky130_fd_sc_hd__o211a_1 _14921_ (.A1(_07621_),
    .A2(_07622_),
    .B1(_07623_),
    .C1(_07620_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _14922_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .S(_07616_),
    .X(_07624_));
 sky130_fd_sc_hd__or2_1 _14923_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(_07618_),
    .X(_07625_));
 sky130_fd_sc_hd__o211a_1 _14924_ (.A1(_07621_),
    .A2(_07624_),
    .B1(_07625_),
    .C1(_07620_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _14925_ (.A0(\rbzero.wall_tracer.trackDistY[0] ),
    .A1(\rbzero.wall_tracer.trackDistX[0] ),
    .S(_07616_),
    .X(_07626_));
 sky130_fd_sc_hd__or2_1 _14926_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .B(_07618_),
    .X(_07627_));
 sky130_fd_sc_hd__o211a_1 _14927_ (.A1(_07621_),
    .A2(_07626_),
    .B1(_07627_),
    .C1(_07620_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _14928_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(\rbzero.wall_tracer.trackDistX[1] ),
    .S(_07616_),
    .X(_07628_));
 sky130_fd_sc_hd__or2_1 _14929_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_07618_),
    .X(_07629_));
 sky130_fd_sc_hd__o211a_1 _14930_ (.A1(_07621_),
    .A2(_07628_),
    .B1(_07629_),
    .C1(_07620_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(\rbzero.wall_tracer.trackDistY[2] ),
    .A1(\rbzero.wall_tracer.trackDistX[2] ),
    .S(_07616_),
    .X(_07630_));
 sky130_fd_sc_hd__or2_1 _14932_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_07618_),
    .X(_07631_));
 sky130_fd_sc_hd__o211a_1 _14933_ (.A1(_07621_),
    .A2(_07630_),
    .B1(_07631_),
    .C1(_07620_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _14934_ (.A0(\rbzero.wall_tracer.trackDistY[3] ),
    .A1(\rbzero.wall_tracer.trackDistX[3] ),
    .S(_07616_),
    .X(_07632_));
 sky130_fd_sc_hd__or2_1 _14935_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_07618_),
    .X(_07633_));
 sky130_fd_sc_hd__o211a_1 _14936_ (.A1(_07621_),
    .A2(_07632_),
    .B1(_07633_),
    .C1(_07620_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _14937_ (.A0(\rbzero.wall_tracer.trackDistY[4] ),
    .A1(\rbzero.wall_tracer.trackDistX[4] ),
    .S(_07616_),
    .X(_07634_));
 sky130_fd_sc_hd__or2_1 _14938_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_07618_),
    .X(_07635_));
 sky130_fd_sc_hd__o211a_1 _14939_ (.A1(_07621_),
    .A2(_07634_),
    .B1(_07635_),
    .C1(_07620_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _14940_ (.A0(\rbzero.wall_tracer.trackDistY[5] ),
    .A1(\rbzero.wall_tracer.trackDistX[5] ),
    .S(_07616_),
    .X(_07636_));
 sky130_fd_sc_hd__or2_1 _14941_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_07618_),
    .X(_07637_));
 sky130_fd_sc_hd__o211a_1 _14942_ (.A1(_07621_),
    .A2(_07636_),
    .B1(_07637_),
    .C1(_07620_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _14943_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(\rbzero.wall_tracer.trackDistX[6] ),
    .S(_07616_),
    .X(_07638_));
 sky130_fd_sc_hd__or2_1 _14944_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_07618_),
    .X(_07639_));
 sky130_fd_sc_hd__o211a_1 _14945_ (.A1(_07621_),
    .A2(_07638_),
    .B1(_07639_),
    .C1(_07620_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _14946_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(\rbzero.wall_tracer.trackDistX[7] ),
    .S(_05278_),
    .X(_07640_));
 sky130_fd_sc_hd__or2_1 _14947_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_07594_),
    .X(_07641_));
 sky130_fd_sc_hd__clkbuf_4 _14948_ (.A(_04035_),
    .X(_07642_));
 sky130_fd_sc_hd__o211a_1 _14949_ (.A1(_07621_),
    .A2(_07640_),
    .B1(_07641_),
    .C1(_07642_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _14950_ (.A0(\rbzero.wall_tracer.trackDistY[8] ),
    .A1(\rbzero.wall_tracer.trackDistX[8] ),
    .S(_05278_),
    .X(_07643_));
 sky130_fd_sc_hd__or2_1 _14951_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_07594_),
    .X(_07644_));
 sky130_fd_sc_hd__o211a_1 _14952_ (.A1(_04019_),
    .A2(_07643_),
    .B1(_07644_),
    .C1(_07642_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _14953_ (.A0(\rbzero.wall_tracer.trackDistY[9] ),
    .A1(\rbzero.wall_tracer.trackDistX[9] ),
    .S(_05278_),
    .X(_07645_));
 sky130_fd_sc_hd__or2_1 _14954_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_07594_),
    .X(_07646_));
 sky130_fd_sc_hd__o211a_1 _14955_ (.A1(_04019_),
    .A2(_07645_),
    .B1(_07646_),
    .C1(_07642_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _14956_ (.A0(\rbzero.wall_tracer.trackDistY[10] ),
    .A1(\rbzero.wall_tracer.trackDistX[10] ),
    .S(_05278_),
    .X(_07647_));
 sky130_fd_sc_hd__or2_1 _14957_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_07594_),
    .X(_07648_));
 sky130_fd_sc_hd__o211a_1 _14958_ (.A1(_04019_),
    .A2(_07647_),
    .B1(_07648_),
    .C1(_07642_),
    .X(_00465_));
 sky130_fd_sc_hd__a21o_1 _14959_ (.A1(\rbzero.wall_tracer.trackDistX[11] ),
    .A2(\rbzero.wall_tracer.trackDistY[11] ),
    .B1(_04019_),
    .X(_07649_));
 sky130_fd_sc_hd__o211a_1 _14960_ (.A1(\rbzero.wall_tracer.visualWallDist[11] ),
    .A2(_07595_),
    .B1(_07649_),
    .C1(_07642_),
    .X(_00466_));
 sky130_fd_sc_hd__buf_4 _14961_ (.A(_05201_),
    .X(_07650_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(\rbzero.wall_tracer.stepDistX[-12] ),
    .A1(_07460_),
    .S(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_07651_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _14964_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_07465_),
    .S(_07650_),
    .X(_07652_));
 sky130_fd_sc_hd__clkbuf_1 _14965_ (.A(_07652_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _14966_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_07484_),
    .S(_07650_),
    .X(_07653_));
 sky130_fd_sc_hd__clkbuf_1 _14967_ (.A(_07653_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _14968_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_07502_),
    .S(_07650_),
    .X(_07654_));
 sky130_fd_sc_hd__clkbuf_1 _14969_ (.A(_07654_),
    .X(_00470_));
 sky130_fd_sc_hd__nor2_1 _14970_ (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .B(_00008_),
    .Y(_07655_));
 sky130_fd_sc_hd__a21oi_1 _14971_ (.A1(_00008_),
    .A2(_07514_),
    .B1(_07655_),
    .Y(_00471_));
 sky130_fd_sc_hd__nor2_1 _14972_ (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .B(_00008_),
    .Y(_07656_));
 sky130_fd_sc_hd__a21oi_1 _14973_ (.A1(_00008_),
    .A2(_07524_),
    .B1(_07656_),
    .Y(_00472_));
 sky130_fd_sc_hd__nor2_1 _14974_ (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .B(_07650_),
    .Y(_07657_));
 sky130_fd_sc_hd__a21oi_1 _14975_ (.A1(_00008_),
    .A2(_07530_),
    .B1(_07657_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2_1 _14976_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_07650_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21oi_1 _14977_ (.A1(_00008_),
    .A2(_07536_),
    .B1(_07658_),
    .Y(_00474_));
 sky130_fd_sc_hd__mux2_1 _14978_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_07541_),
    .S(_07650_),
    .X(_07659_));
 sky130_fd_sc_hd__clkbuf_1 _14979_ (.A(_07659_),
    .X(_00475_));
 sky130_fd_sc_hd__buf_4 _14980_ (.A(_05201_),
    .X(_07660_));
 sky130_fd_sc_hd__mux2_1 _14981_ (.A0(\rbzero.wall_tracer.stepDistX[-3] ),
    .A1(_07545_),
    .S(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__clkbuf_1 _14982_ (.A(_07661_),
    .X(_00476_));
 sky130_fd_sc_hd__nor2_1 _14983_ (.A(\rbzero.wall_tracer.stepDistX[-2] ),
    .B(_07650_),
    .Y(_07662_));
 sky130_fd_sc_hd__a21oi_1 _14984_ (.A1(_00008_),
    .A2(_07549_),
    .B1(_07662_),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_1 _14985_ (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .B(_07650_),
    .Y(_07663_));
 sky130_fd_sc_hd__a21oi_1 _14986_ (.A1(_00008_),
    .A2(_07552_),
    .B1(_07663_),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_1 _14987_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .B(_07650_),
    .Y(_07664_));
 sky130_fd_sc_hd__a21oi_1 _14988_ (.A1(_00008_),
    .A2(_07555_),
    .B1(_07664_),
    .Y(_00479_));
 sky130_fd_sc_hd__mux2_1 _14989_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_07560_),
    .S(_07660_),
    .X(_07665_));
 sky130_fd_sc_hd__clkbuf_1 _14990_ (.A(_07665_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _14991_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_07562_),
    .S(_07660_),
    .X(_07666_));
 sky130_fd_sc_hd__clkbuf_1 _14992_ (.A(_07666_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _14993_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_07564_),
    .S(_07660_),
    .X(_07667_));
 sky130_fd_sc_hd__clkbuf_1 _14994_ (.A(_07667_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _14995_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_07566_),
    .S(_07660_),
    .X(_07668_));
 sky130_fd_sc_hd__clkbuf_1 _14996_ (.A(_07668_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _14997_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_07568_),
    .S(_07660_),
    .X(_07669_));
 sky130_fd_sc_hd__clkbuf_1 _14998_ (.A(_07669_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _14999_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_07571_),
    .S(_07660_),
    .X(_07670_));
 sky130_fd_sc_hd__clkbuf_1 _15000_ (.A(_07670_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _15001_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_07575_),
    .S(_07660_),
    .X(_07671_));
 sky130_fd_sc_hd__clkbuf_1 _15002_ (.A(_07671_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _15003_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_07579_),
    .S(_07660_),
    .X(_07672_));
 sky130_fd_sc_hd__clkbuf_1 _15004_ (.A(_07672_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _15005_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_07582_),
    .S(_07660_),
    .X(_07673_));
 sky130_fd_sc_hd__clkbuf_1 _15006_ (.A(_07673_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _15007_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_07586_),
    .S(_05201_),
    .X(_07674_));
 sky130_fd_sc_hd__clkbuf_1 _15008_ (.A(_07674_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _15009_ (.A0(\rbzero.wall_tracer.stepDistX[11] ),
    .A1(_07589_),
    .S(_05201_),
    .X(_07675_));
 sky130_fd_sc_hd__clkbuf_1 _15010_ (.A(_07675_),
    .X(_00490_));
 sky130_fd_sc_hd__clkbuf_4 _15011_ (.A(_03912_),
    .X(_07676_));
 sky130_fd_sc_hd__nand2_2 _15012_ (.A(\rbzero.wall_tracer.state[14] ),
    .B(_04037_),
    .Y(_07677_));
 sky130_fd_sc_hd__nor2_1 _15013_ (.A(_07676_),
    .B(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__buf_4 _15014_ (.A(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__nor2_1 _15015_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_07680_));
 sky130_fd_sc_hd__nand2_1 _15016_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_07681_));
 sky130_fd_sc_hd__and2b_1 _15017_ (.A_N(_07680_),
    .B(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__or2_1 _15018_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .X(_07683_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_07684_));
 sky130_fd_sc_hd__nand2_1 _15020_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .Y(_07685_));
 sky130_fd_sc_hd__or2_1 _15021_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_07686_));
 sky130_fd_sc_hd__nand2_1 _15022_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_07687_));
 sky130_fd_sc_hd__and3b_1 _15023_ (.A_N(_07685_),
    .B(_07686_),
    .C(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__a21oi_1 _15024_ (.A1(\rbzero.debug_overlay.vplaneX[-8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-8] ),
    .B1(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__nand2_1 _15025_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_07690_));
 sky130_fd_sc_hd__o21ai_2 _15026_ (.A1(_07684_),
    .A2(_07689_),
    .B1(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_07692_));
 sky130_fd_sc_hd__a21boi_1 _15028_ (.A1(_07683_),
    .A2(_07691_),
    .B1_N(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__xnor2_1 _15029_ (.A(_07682_),
    .B(_07693_),
    .Y(_07694_));
 sky130_fd_sc_hd__buf_4 _15030_ (.A(_04028_),
    .X(_07695_));
 sky130_fd_sc_hd__and2_1 _15031_ (.A(\rbzero.wall_tracer.rayAddendX[-5] ),
    .B(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__a221o_1 _15032_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_03914_),
    .B1(_07679_),
    .B2(_07694_),
    .C1(_07696_),
    .X(_00491_));
 sky130_fd_sc_hd__nor2_1 _15033_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_07697_));
 sky130_fd_sc_hd__and2_1 _15034_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_07698_));
 sky130_fd_sc_hd__o21ai_1 _15035_ (.A1(_07680_),
    .A2(_07693_),
    .B1(_07681_),
    .Y(_07699_));
 sky130_fd_sc_hd__or3_1 _15036_ (.A(_07697_),
    .B(_07698_),
    .C(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__o21ai_1 _15037_ (.A1(_07697_),
    .A2(_07698_),
    .B1(_07699_),
    .Y(_07701_));
 sky130_fd_sc_hd__a21oi_1 _15038_ (.A1(_07700_),
    .A2(_07701_),
    .B1(_03914_),
    .Y(_07702_));
 sky130_fd_sc_hd__clkbuf_4 _15039_ (.A(_03913_),
    .X(_07703_));
 sky130_fd_sc_hd__nand2_1 _15040_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_07704_));
 sky130_fd_sc_hd__or2_1 _15041_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_07705_));
 sky130_fd_sc_hd__buf_4 _15042_ (.A(_07695_),
    .X(_07706_));
 sky130_fd_sc_hd__a31o_1 _15043_ (.A1(_07703_),
    .A2(_07704_),
    .A3(_07705_),
    .B1(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__o22a_1 _15044_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_00013_),
    .B1(_07702_),
    .B2(_07707_),
    .X(_00492_));
 sky130_fd_sc_hd__or2_1 _15045_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_07705_),
    .X(_07708_));
 sky130_fd_sc_hd__nand2_1 _15046_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_07705_),
    .Y(_07709_));
 sky130_fd_sc_hd__nor2_1 _15047_ (.A(_04462_),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_07710_));
 sky130_fd_sc_hd__nand2_1 _15048_ (.A(_04462_),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_07711_));
 sky130_fd_sc_hd__or2b_1 _15049_ (.A(_07710_),
    .B_N(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__or2_1 _15050_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_07713_));
 sky130_fd_sc_hd__a21oi_1 _15051_ (.A1(_07713_),
    .A2(_07699_),
    .B1(_07698_),
    .Y(_07714_));
 sky130_fd_sc_hd__xnor2_1 _15052_ (.A(_07712_),
    .B(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__nor2_1 _15053_ (.A(_07676_),
    .B(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__a31o_1 _15054_ (.A1(_07676_),
    .A2(_07708_),
    .A3(_07709_),
    .B1(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__buf_4 _15055_ (.A(_04029_),
    .X(_07718_));
 sky130_fd_sc_hd__mux2_1 _15056_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_07717_),
    .S(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__clkbuf_1 _15057_ (.A(_07719_),
    .X(_00493_));
 sky130_fd_sc_hd__xor2_1 _15058_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_07708_),
    .X(_07720_));
 sky130_fd_sc_hd__or2_1 _15059_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_07721_));
 sky130_fd_sc_hd__nand2_1 _15060_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_07722_));
 sky130_fd_sc_hd__nand2_1 _15061_ (.A(_07721_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__o21ai_1 _15062_ (.A1(_07710_),
    .A2(_07714_),
    .B1(_07711_),
    .Y(_07724_));
 sky130_fd_sc_hd__xnor2_1 _15063_ (.A(_07723_),
    .B(_07724_),
    .Y(_07725_));
 sky130_fd_sc_hd__mux2_1 _15064_ (.A0(_07720_),
    .A1(_07725_),
    .S(_04033_),
    .X(_07726_));
 sky130_fd_sc_hd__mux2_1 _15065_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_07726_),
    .S(_07718_),
    .X(_07727_));
 sky130_fd_sc_hd__clkbuf_1 _15066_ (.A(_07727_),
    .X(_00494_));
 sky130_fd_sc_hd__buf_4 _15067_ (.A(_07679_),
    .X(_07728_));
 sky130_fd_sc_hd__or2_1 _15068_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_07729_));
 sky130_fd_sc_hd__clkbuf_4 _15069_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_07730_));
 sky130_fd_sc_hd__nand2_1 _15070_ (.A(_07730_),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_07731_));
 sky130_fd_sc_hd__nand2_1 _15071_ (.A(_07729_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__a21bo_1 _15072_ (.A1(_07721_),
    .A2(_07724_),
    .B1_N(_07722_),
    .X(_07733_));
 sky130_fd_sc_hd__xnor2_1 _15073_ (.A(_07732_),
    .B(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__or4b_1 _15074_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .C(\rbzero.debug_overlay.vplaneX[-9] ),
    .D_N(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_07735_));
 sky130_fd_sc_hd__or2_1 _15075_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_07736_));
 sky130_fd_sc_hd__nand2_1 _15076_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_07737_));
 sky130_fd_sc_hd__a2bb2o_1 _15077_ (.A1_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2_N(_07708_),
    .B1(_07736_),
    .B2(_07737_),
    .X(_07738_));
 sky130_fd_sc_hd__o21ai_1 _15078_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(_07735_),
    .B1(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__a22o_1 _15079_ (.A1(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2(_07706_),
    .B1(_07739_),
    .B2(_07703_),
    .X(_07740_));
 sky130_fd_sc_hd__a21o_1 _15080_ (.A1(_07728_),
    .A2(_07734_),
    .B1(_07740_),
    .X(_00495_));
 sky130_fd_sc_hd__a21bo_1 _15081_ (.A1(_07729_),
    .A2(_07733_),
    .B1_N(_07731_),
    .X(_07741_));
 sky130_fd_sc_hd__buf_2 _15082_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_07742_));
 sky130_fd_sc_hd__nor2_1 _15083_ (.A(_07742_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_07743_));
 sky130_fd_sc_hd__and2_1 _15084_ (.A(_07742_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_07744_));
 sky130_fd_sc_hd__nor2_1 _15085_ (.A(_07743_),
    .B(_07744_),
    .Y(_07745_));
 sky130_fd_sc_hd__o21ai_1 _15086_ (.A1(_07741_),
    .A2(_07745_),
    .B1(_04034_),
    .Y(_07746_));
 sky130_fd_sc_hd__a21oi_1 _15087_ (.A1(_07741_),
    .A2(_07745_),
    .B1(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__and2_1 _15088_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_07748_));
 sky130_fd_sc_hd__nor2_1 _15089_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .Y(_07749_));
 sky130_fd_sc_hd__o21ai_1 _15090_ (.A1(_07748_),
    .A2(_07749_),
    .B1(_07736_),
    .Y(_07750_));
 sky130_fd_sc_hd__or3_1 _15091_ (.A(_07736_),
    .B(_07748_),
    .C(_07749_),
    .X(_07751_));
 sky130_fd_sc_hd__and2_1 _15092_ (.A(_07750_),
    .B(_07751_),
    .X(_07752_));
 sky130_fd_sc_hd__or2_1 _15093_ (.A(_07738_),
    .B(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__nand2_1 _15094_ (.A(_07738_),
    .B(_07752_),
    .Y(_07754_));
 sky130_fd_sc_hd__a31o_1 _15095_ (.A1(_07703_),
    .A2(_07753_),
    .A3(_07754_),
    .B1(_07706_),
    .X(_07755_));
 sky130_fd_sc_hd__o22a_1 _15096_ (.A1(\rbzero.wall_tracer.rayAddendX[0] ),
    .A2(_00013_),
    .B1(_07747_),
    .B2(_07755_),
    .X(_00496_));
 sky130_fd_sc_hd__buf_6 _15097_ (.A(_07678_),
    .X(_07756_));
 sky130_fd_sc_hd__or2_1 _15098_ (.A(_07742_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_07757_));
 sky130_fd_sc_hd__nand2_1 _15099_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_07758_));
 sky130_fd_sc_hd__or2_1 _15100_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_07759_));
 sky130_fd_sc_hd__or2_1 _15101_ (.A(_07741_),
    .B(_07744_),
    .X(_07760_));
 sky130_fd_sc_hd__nand4_2 _15102_ (.A(_07757_),
    .B(_07758_),
    .C(_07759_),
    .D(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__a22o_1 _15103_ (.A1(_07758_),
    .A2(_07759_),
    .B1(_07760_),
    .B2(_07757_),
    .X(_07762_));
 sky130_fd_sc_hd__xnor2_1 _15104_ (.A(_04462_),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_07763_));
 sky130_fd_sc_hd__a21oi_1 _15105_ (.A1(_07751_),
    .A2(_07754_),
    .B1(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__and3_1 _15106_ (.A(_07751_),
    .B(_07754_),
    .C(_07763_),
    .X(_07765_));
 sky130_fd_sc_hd__or2_1 _15107_ (.A(_07764_),
    .B(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__xnor2_1 _15108_ (.A(_07749_),
    .B(_07766_),
    .Y(_07767_));
 sky130_fd_sc_hd__a22o_1 _15109_ (.A1(\rbzero.wall_tracer.rayAddendX[1] ),
    .A2(_07695_),
    .B1(_07767_),
    .B2(_07703_),
    .X(_07768_));
 sky130_fd_sc_hd__a31o_1 _15110_ (.A1(_07756_),
    .A2(_07761_),
    .A3(_07762_),
    .B1(_07768_),
    .X(_00497_));
 sky130_fd_sc_hd__nand2_1 _15111_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_07769_));
 sky130_fd_sc_hd__or2_1 _15112_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .X(_07770_));
 sky130_fd_sc_hd__nand2_1 _15113_ (.A(_07769_),
    .B(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__a21oi_1 _15114_ (.A1(_07758_),
    .A2(_07761_),
    .B1(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__a31o_1 _15115_ (.A1(_07758_),
    .A2(_07761_),
    .A3(_07771_),
    .B1(_03912_),
    .X(_07773_));
 sky130_fd_sc_hd__and2_1 _15116_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_07774_));
 sky130_fd_sc_hd__nor2_1 _15117_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .Y(_07775_));
 sky130_fd_sc_hd__o22a_1 _15118_ (.A1(_04462_),
    .A2(\rbzero.debug_overlay.vplaneX[-7] ),
    .B1(_07774_),
    .B2(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__nor4_1 _15119_ (.A(_04462_),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .C(_07774_),
    .D(_07775_),
    .Y(_07777_));
 sky130_fd_sc_hd__or2_1 _15120_ (.A(_07776_),
    .B(_07777_),
    .X(_07778_));
 sky130_fd_sc_hd__o2bb2ai_1 _15121_ (.A1_N(_07754_),
    .A2_N(_07763_),
    .B1(_07764_),
    .B2(_07749_),
    .Y(_07779_));
 sky130_fd_sc_hd__xor2_1 _15122_ (.A(_07778_),
    .B(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__a2bb2o_1 _15123_ (.A1_N(_07772_),
    .A2_N(_07773_),
    .B1(_07780_),
    .B2(_07676_),
    .X(_07781_));
 sky130_fd_sc_hd__mux2_1 _15124_ (.A0(\rbzero.wall_tracer.rayAddendX[2] ),
    .A1(_07781_),
    .S(_07718_),
    .X(_07782_));
 sky130_fd_sc_hd__clkbuf_1 _15125_ (.A(_07782_),
    .X(_00498_));
 sky130_fd_sc_hd__nor2_1 _15126_ (.A(_07761_),
    .B(_07771_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand2_1 _15127_ (.A(_07758_),
    .B(_07769_),
    .Y(_07784_));
 sky130_fd_sc_hd__clkbuf_4 _15128_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_07785_));
 sky130_fd_sc_hd__nand2_1 _15129_ (.A(_07785_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_07786_));
 sky130_fd_sc_hd__or2_1 _15130_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_07787_));
 sky130_fd_sc_hd__o211a_1 _15131_ (.A1(_07783_),
    .A2(_07784_),
    .B1(_07786_),
    .C1(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__inv_2 _15132_ (.A(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__a211o_1 _15133_ (.A1(_07786_),
    .A2(_07787_),
    .B1(_07783_),
    .C1(_07784_),
    .X(_07790_));
 sky130_fd_sc_hd__xor2_1 _15134_ (.A(_07730_),
    .B(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_07791_));
 sky130_fd_sc_hd__nor2_1 _15135_ (.A(_07778_),
    .B(_07779_),
    .Y(_07792_));
 sky130_fd_sc_hd__or2_1 _15136_ (.A(_07777_),
    .B(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__xnor2_1 _15137_ (.A(_07791_),
    .B(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__xnor2_1 _15138_ (.A(_07775_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__a22o_1 _15139_ (.A1(\rbzero.wall_tracer.rayAddendX[3] ),
    .A2(_07695_),
    .B1(_07795_),
    .B2(_07703_),
    .X(_07796_));
 sky130_fd_sc_hd__a31o_1 _15140_ (.A1(_07756_),
    .A2(_07789_),
    .A3(_07790_),
    .B1(_07796_),
    .X(_00499_));
 sky130_fd_sc_hd__xor2_1 _15141_ (.A(_07785_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_07797_));
 sky130_fd_sc_hd__and2_1 _15142_ (.A(_07786_),
    .B(_07789_),
    .X(_07798_));
 sky130_fd_sc_hd__xnor2_1 _15143_ (.A(_07797_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__nor2_1 _15144_ (.A(_07742_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .Y(_07800_));
 sky130_fd_sc_hd__and2_1 _15145_ (.A(_07742_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_07801_));
 sky130_fd_sc_hd__o22a_1 _15146_ (.A1(_07730_),
    .A2(\rbzero.debug_overlay.vplaneX[-5] ),
    .B1(_07800_),
    .B2(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__nor4_1 _15147_ (.A(_07730_),
    .B(\rbzero.debug_overlay.vplaneX[-5] ),
    .C(_07800_),
    .D(_07801_),
    .Y(_07803_));
 sky130_fd_sc_hd__nor2_1 _15148_ (.A(_07802_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__and2_1 _15149_ (.A(_07791_),
    .B(_07793_),
    .X(_07805_));
 sky130_fd_sc_hd__o22a_1 _15150_ (.A1(_07792_),
    .A2(_07791_),
    .B1(_07805_),
    .B2(_07775_),
    .X(_07806_));
 sky130_fd_sc_hd__or2_1 _15151_ (.A(_07804_),
    .B(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__and2_1 _15152_ (.A(_07804_),
    .B(_07806_),
    .X(_07808_));
 sky130_fd_sc_hd__nor2_1 _15153_ (.A(_04033_),
    .B(_07808_),
    .Y(_07809_));
 sky130_fd_sc_hd__a22o_1 _15154_ (.A1(_04034_),
    .A2(_07799_),
    .B1(_07807_),
    .B2(_07809_),
    .X(_07810_));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_07810_),
    .S(_07718_),
    .X(_07811_));
 sky130_fd_sc_hd__clkbuf_1 _15156_ (.A(_07811_),
    .X(_00500_));
 sky130_fd_sc_hd__xor2_1 _15157_ (.A(_07785_),
    .B(_04462_),
    .X(_07812_));
 sky130_fd_sc_hd__xor2_1 _15158_ (.A(_07800_),
    .B(_07812_),
    .X(_07813_));
 sky130_fd_sc_hd__o21a_1 _15159_ (.A1(_07803_),
    .A2(_07808_),
    .B1(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__o31ai_1 _15160_ (.A1(_07803_),
    .A2(_07808_),
    .A3(_07813_),
    .B1(_07676_),
    .Y(_07815_));
 sky130_fd_sc_hd__nand2_1 _15161_ (.A(_07785_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_07816_));
 sky130_fd_sc_hd__or2_1 _15162_ (.A(_07785_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_07817_));
 sky130_fd_sc_hd__nand2_1 _15163_ (.A(_07816_),
    .B(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__nand2_1 _15164_ (.A(_07788_),
    .B(_07797_),
    .Y(_07819_));
 sky130_fd_sc_hd__buf_2 _15165_ (.A(_07785_),
    .X(_07820_));
 sky130_fd_sc_hd__clkbuf_4 _15166_ (.A(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__o21ai_1 _15167_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__and3_1 _15168_ (.A(_07818_),
    .B(_07819_),
    .C(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__a21o_1 _15169_ (.A1(_07819_),
    .A2(_07822_),
    .B1(_07818_),
    .X(_07824_));
 sky130_fd_sc_hd__and2b_1 _15170_ (.A_N(_07823_),
    .B(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__a2bb2o_1 _15171_ (.A1_N(_07814_),
    .A2_N(_07815_),
    .B1(_04033_),
    .B2(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__mux2_1 _15172_ (.A0(\rbzero.wall_tracer.rayAddendX[5] ),
    .A1(_07826_),
    .S(_07718_),
    .X(_07827_));
 sky130_fd_sc_hd__clkbuf_1 _15173_ (.A(_07827_),
    .X(_00501_));
 sky130_fd_sc_hd__xnor2_1 _15174_ (.A(_07785_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_07828_));
 sky130_fd_sc_hd__a21oi_1 _15175_ (.A1(_07816_),
    .A2(_07824_),
    .B1(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand2_8 _15176_ (.A(_04033_),
    .B(_04027_),
    .Y(_07830_));
 sky130_fd_sc_hd__buf_6 _15177_ (.A(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__a31o_1 _15178_ (.A1(_07816_),
    .A2(_07824_),
    .A3(_07828_),
    .B1(_07831_),
    .X(_07832_));
 sky130_fd_sc_hd__nor2_1 _15179_ (.A(_07820_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .Y(_07833_));
 sky130_fd_sc_hd__and2_1 _15180_ (.A(_07785_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_07834_));
 sky130_fd_sc_hd__o22ai_1 _15181_ (.A1(_07820_),
    .A2(_04462_),
    .B1(_07833_),
    .B2(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__or3b_1 _15182_ (.A(_07820_),
    .B(_04462_),
    .C_N(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_07836_));
 sky130_fd_sc_hd__nand2_1 _15183_ (.A(_07835_),
    .B(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__a21o_1 _15184_ (.A1(_07800_),
    .A2(_07812_),
    .B1(_07814_),
    .X(_07838_));
 sky130_fd_sc_hd__xnor2_1 _15185_ (.A(_07837_),
    .B(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__a22o_1 _15186_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_07695_),
    .B1(_07839_),
    .B2(_03913_),
    .X(_07840_));
 sky130_fd_sc_hd__o21bai_1 _15187_ (.A1(_07829_),
    .A2(_07832_),
    .B1_N(_07840_),
    .Y(_00502_));
 sky130_fd_sc_hd__nor3_1 _15188_ (.A(_07818_),
    .B(_07819_),
    .C(_07828_),
    .Y(_07841_));
 sky130_fd_sc_hd__o41a_1 _15189_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .A3(\rbzero.wall_tracer.rayAddendX[4] ),
    .A4(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_07785_),
    .X(_07842_));
 sky130_fd_sc_hd__nand2_1 _15190_ (.A(_07820_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_07843_));
 sky130_fd_sc_hd__or2_1 _15191_ (.A(_07785_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_07844_));
 sky130_fd_sc_hd__o211ai_2 _15192_ (.A1(_07841_),
    .A2(_07842_),
    .B1(_07843_),
    .C1(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__a211o_1 _15193_ (.A1(_07843_),
    .A2(_07844_),
    .B1(_07841_),
    .C1(_07842_),
    .X(_07846_));
 sky130_fd_sc_hd__nor2_1 _15194_ (.A(_07820_),
    .B(_07730_),
    .Y(_07847_));
 sky130_fd_sc_hd__and2_1 _15195_ (.A(_07820_),
    .B(_07730_),
    .X(_07848_));
 sky130_fd_sc_hd__o21bai_1 _15196_ (.A1(_07847_),
    .A2(_07848_),
    .B1_N(_07833_),
    .Y(_07849_));
 sky130_fd_sc_hd__nand2_1 _15197_ (.A(_07730_),
    .B(_07833_),
    .Y(_07850_));
 sky130_fd_sc_hd__nand2_1 _15198_ (.A(_07849_),
    .B(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__a21boi_1 _15199_ (.A1(_07835_),
    .A2(_07838_),
    .B1_N(_07836_),
    .Y(_07852_));
 sky130_fd_sc_hd__nand2_1 _15200_ (.A(_07851_),
    .B(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__or2_1 _15201_ (.A(_07851_),
    .B(_07852_),
    .X(_07854_));
 sky130_fd_sc_hd__buf_4 _15202_ (.A(_04028_),
    .X(_07855_));
 sky130_fd_sc_hd__a32o_1 _15203_ (.A1(_03913_),
    .A2(_07853_),
    .A3(_07854_),
    .B1(_07855_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_07856_));
 sky130_fd_sc_hd__a31o_1 _15204_ (.A1(_07756_),
    .A2(_07845_),
    .A3(_07846_),
    .B1(_07856_),
    .X(_00503_));
 sky130_fd_sc_hd__nand2_1 _15205_ (.A(_07821_),
    .B(_07742_),
    .Y(_07857_));
 sky130_fd_sc_hd__or2_1 _15206_ (.A(_07821_),
    .B(_07742_),
    .X(_07858_));
 sky130_fd_sc_hd__a21oi_1 _15207_ (.A1(_07857_),
    .A2(_07858_),
    .B1(_07847_),
    .Y(_07859_));
 sky130_fd_sc_hd__a21o_1 _15208_ (.A1(_07742_),
    .A2(_07847_),
    .B1(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__and3_1 _15209_ (.A(_07850_),
    .B(_07854_),
    .C(_07860_),
    .X(_07861_));
 sky130_fd_sc_hd__a21oi_1 _15210_ (.A1(_07850_),
    .A2(_07854_),
    .B1(_07860_),
    .Y(_07862_));
 sky130_fd_sc_hd__o31a_1 _15211_ (.A1(_04034_),
    .A2(_07861_),
    .A3(_07862_),
    .B1(_07718_),
    .X(_07863_));
 sky130_fd_sc_hd__xnor2_1 _15212_ (.A(_07820_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_07864_));
 sky130_fd_sc_hd__a21oi_1 _15213_ (.A1(_07843_),
    .A2(_07845_),
    .B1(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__a31o_1 _15214_ (.A1(_07843_),
    .A2(_07845_),
    .A3(_07864_),
    .B1(_07676_),
    .X(_07866_));
 sky130_fd_sc_hd__or2_1 _15215_ (.A(_07865_),
    .B(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__o2bb2a_1 _15216_ (.A1_N(_07863_),
    .A2_N(_07867_),
    .B1(_00013_),
    .B2(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_00504_));
 sky130_fd_sc_hd__nor2_1 _15217_ (.A(_07845_),
    .B(_07864_),
    .Y(_07868_));
 sky130_fd_sc_hd__o21a_1 _15218_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .B1(_07821_),
    .X(_07869_));
 sky130_fd_sc_hd__nand2_1 _15219_ (.A(_07820_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_07870_));
 sky130_fd_sc_hd__or2_1 _15220_ (.A(_07820_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_07871_));
 sky130_fd_sc_hd__and2_1 _15221_ (.A(_07870_),
    .B(_07871_),
    .X(_07872_));
 sky130_fd_sc_hd__o21ai_1 _15222_ (.A1(_07868_),
    .A2(_07869_),
    .B1(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__or3_1 _15223_ (.A(_07872_),
    .B(_07868_),
    .C(_07869_),
    .X(_07874_));
 sky130_fd_sc_hd__and2_1 _15224_ (.A(_07873_),
    .B(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__a211oi_1 _15225_ (.A1(_07742_),
    .A2(_07730_),
    .B1(_07862_),
    .C1(_07821_),
    .Y(_07876_));
 sky130_fd_sc_hd__a211o_1 _15226_ (.A1(_07858_),
    .A2(_07862_),
    .B1(_07876_),
    .C1(_04034_),
    .X(_07877_));
 sky130_fd_sc_hd__o221a_1 _15227_ (.A1(\rbzero.wall_tracer.rayAddendX[9] ),
    .A2(_00013_),
    .B1(_07831_),
    .B2(_07875_),
    .C1(_07877_),
    .X(_00505_));
 sky130_fd_sc_hd__nor2_1 _15228_ (.A(_07730_),
    .B(_07854_),
    .Y(_07878_));
 sky130_fd_sc_hd__or3_1 _15229_ (.A(_07821_),
    .B(_04033_),
    .C(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__inv_2 _15230_ (.A(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__xnor2_1 _15231_ (.A(_07821_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_07881_));
 sky130_fd_sc_hd__a21oi_1 _15232_ (.A1(_07870_),
    .A2(_07873_),
    .B1(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__a31o_1 _15233_ (.A1(_07870_),
    .A2(_07873_),
    .A3(_07881_),
    .B1(_07830_),
    .X(_07883_));
 sky130_fd_sc_hd__nor2_1 _15234_ (.A(_07882_),
    .B(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__a211o_1 _15235_ (.A1(\rbzero.wall_tracer.rayAddendX[10] ),
    .A2(_07855_),
    .B1(_07880_),
    .C1(_07884_),
    .X(_00506_));
 sky130_fd_sc_hd__or4b_1 _15236_ (.A(\rbzero.wall_tracer.rayAddendX[8] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .C(_05448_),
    .D_N(_07821_),
    .X(_07885_));
 sky130_fd_sc_hd__and3b_1 _15237_ (.A_N(_07881_),
    .B(_07868_),
    .C(_07872_),
    .X(_07886_));
 sky130_fd_sc_hd__mux2_1 _15238_ (.A0(_07885_),
    .A1(_07821_),
    .S(_07886_),
    .X(_07887_));
 sky130_fd_sc_hd__xnor2_1 _15239_ (.A(\rbzero.wall_tracer.rayAddendX[11] ),
    .B(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__a221o_1 _15240_ (.A1(\rbzero.wall_tracer.rayAddendX[11] ),
    .A2(_07855_),
    .B1(_07679_),
    .B2(_07888_),
    .C1(_07880_),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _15241_ (.A1(\rbzero.wall_tracer.wall[0] ),
    .A2(_03999_),
    .B1(_05280_),
    .B2(_03987_),
    .X(_07889_));
 sky130_fd_sc_hd__and2_1 _15242_ (.A(_04035_),
    .B(_07889_),
    .X(_07890_));
 sky130_fd_sc_hd__clkbuf_1 _15243_ (.A(_07890_),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _15244_ (.A1(\rbzero.wall_tracer.wall[1] ),
    .A2(_03999_),
    .B1(_05280_),
    .B2(_03996_),
    .X(_07891_));
 sky130_fd_sc_hd__and2_1 _15245_ (.A(_04035_),
    .B(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__clkbuf_1 _15246_ (.A(_07892_),
    .X(_00509_));
 sky130_fd_sc_hd__clkbuf_4 _15247_ (.A(\rbzero.wall_tracer.side ),
    .X(_07893_));
 sky130_fd_sc_hd__clkbuf_4 _15248_ (.A(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__buf_4 _15249_ (.A(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__nand2_1 _15250_ (.A(_07595_),
    .B(_07592_),
    .Y(_07896_));
 sky130_fd_sc_hd__o211a_1 _15251_ (.A1(_07895_),
    .A2(_07595_),
    .B1(_07896_),
    .C1(_07642_),
    .X(_00510_));
 sky130_fd_sc_hd__or3_1 _15252_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_07897_));
 sky130_fd_sc_hd__or2_2 _15253_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__nand2_1 _15254_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_07897_),
    .Y(_07899_));
 sky130_fd_sc_hd__nand2_1 _15255_ (.A(_07898_),
    .B(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__inv_2 _15256_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .Y(_07901_));
 sky130_fd_sc_hd__mux2_1 _15257_ (.A0(_07900_),
    .A1(_07901_),
    .S(_05495_),
    .X(_07902_));
 sky130_fd_sc_hd__clkbuf_4 _15258_ (.A(\rbzero.wall_tracer.state[13] ),
    .X(_07903_));
 sky130_fd_sc_hd__clkbuf_4 _15259_ (.A(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__or3_1 _15260_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_07905_));
 sky130_fd_sc_hd__or2_1 _15261_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__nand2_1 _15262_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_07905_),
    .Y(_07907_));
 sky130_fd_sc_hd__and2_1 _15263_ (.A(_07906_),
    .B(_07907_),
    .X(_07908_));
 sky130_fd_sc_hd__mux2_1 _15264_ (.A0(_07908_),
    .A1(\rbzero.debug_overlay.playerY[-6] ),
    .S(_05373_),
    .X(_07909_));
 sky130_fd_sc_hd__nand2_1 _15265_ (.A(_07904_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__a21oi_1 _15266_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_04013_),
    .B1(_05195_),
    .Y(_07911_));
 sky130_fd_sc_hd__a22o_4 _15267_ (.A1(_05206_),
    .A2(_07902_),
    .B1(_07910_),
    .B2(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__clkbuf_4 _15268_ (.A(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__xnor2_2 _15269_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_07898_),
    .Y(_07914_));
 sky130_fd_sc_hd__nand2_1 _15270_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_05495_),
    .Y(_07915_));
 sky130_fd_sc_hd__o211a_4 _15271_ (.A1(_05495_),
    .A2(_07914_),
    .B1(_07915_),
    .C1(_05195_),
    .X(_07916_));
 sky130_fd_sc_hd__xor2_1 _15272_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_07906_),
    .X(_07917_));
 sky130_fd_sc_hd__mux2_2 _15273_ (.A0(_07917_),
    .A1(\rbzero.debug_overlay.playerY[-5] ),
    .S(_05373_),
    .X(_07918_));
 sky130_fd_sc_hd__a21o_1 _15274_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_04012_),
    .B1(\rbzero.wall_tracer.state[6] ),
    .X(_07919_));
 sky130_fd_sc_hd__a21o_1 _15275_ (.A1(_07903_),
    .A2(_07918_),
    .B1(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__clkinv_2 _15276_ (.A(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__or2_1 _15277_ (.A(_07916_),
    .B(_07921_),
    .X(_07922_));
 sky130_fd_sc_hd__clkbuf_2 _15278_ (.A(_07922_),
    .X(_07923_));
 sky130_fd_sc_hd__buf_2 _15279_ (.A(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__clkbuf_8 _15280_ (.A(_04013_),
    .X(_07925_));
 sky130_fd_sc_hd__mux2_1 _15281_ (.A0(_05346_),
    .A1(_05468_),
    .S(_07893_),
    .X(_07926_));
 sky130_fd_sc_hd__mux2_1 _15282_ (.A0(_07541_),
    .A1(_07926_),
    .S(\rbzero.wall_tracer.state[3] ),
    .X(_07927_));
 sky130_fd_sc_hd__a21o_1 _15283_ (.A1(_07904_),
    .A2(\rbzero.wall_tracer.stepDistY[-4] ),
    .B1(_05195_),
    .X(_07928_));
 sky130_fd_sc_hd__a21oi_1 _15284_ (.A1(_07925_),
    .A2(_07927_),
    .B1(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__nor2_1 _15285_ (.A(_05197_),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_07930_));
 sky130_fd_sc_hd__or2_2 _15286_ (.A(_07929_),
    .B(_07930_),
    .X(_07931_));
 sky130_fd_sc_hd__clkbuf_4 _15287_ (.A(_07931_),
    .X(_07932_));
 sky130_fd_sc_hd__buf_4 _15288_ (.A(\rbzero.wall_tracer.state[3] ),
    .X(_07933_));
 sky130_fd_sc_hd__mux2_1 _15289_ (.A0(_05349_),
    .A1(_05469_),
    .S(\rbzero.wall_tracer.side ),
    .X(_07934_));
 sky130_fd_sc_hd__nand2_1 _15290_ (.A(_07933_),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__o21ai_4 _15291_ (.A1(_07933_),
    .A2(_07536_),
    .B1(_07935_),
    .Y(_07936_));
 sky130_fd_sc_hd__a21o_1 _15292_ (.A1(_07903_),
    .A2(\rbzero.wall_tracer.stepDistY[-5] ),
    .B1(_05195_),
    .X(_07937_));
 sky130_fd_sc_hd__a21oi_4 _15293_ (.A1(_04013_),
    .A2(_07936_),
    .B1(_07937_),
    .Y(_07938_));
 sky130_fd_sc_hd__nor2_2 _15294_ (.A(_05197_),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_07939_));
 sky130_fd_sc_hd__or2_1 _15295_ (.A(_07938_),
    .B(_07939_),
    .X(_07940_));
 sky130_fd_sc_hd__clkbuf_4 _15296_ (.A(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__or4_1 _15297_ (.A(_07913_),
    .B(_07924_),
    .C(_07932_),
    .D(_07941_),
    .X(_07942_));
 sky130_fd_sc_hd__o22ai_1 _15298_ (.A1(_07913_),
    .A2(_07932_),
    .B1(_07941_),
    .B2(_07924_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_1 _15299_ (.A(_07942_),
    .B(_07943_),
    .Y(_07944_));
 sky130_fd_sc_hd__buf_6 _15300_ (.A(_05207_),
    .X(_07945_));
 sky130_fd_sc_hd__or3_1 _15301_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_07898_),
    .X(_07946_));
 sky130_fd_sc_hd__o21ai_1 _15302_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_07898_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_07947_));
 sky130_fd_sc_hd__nand2_1 _15303_ (.A(_07946_),
    .B(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__inv_2 _15304_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_07949_));
 sky130_fd_sc_hd__mux2_1 _15305_ (.A0(_07948_),
    .A1(_07949_),
    .S(_05496_),
    .X(_07950_));
 sky130_fd_sc_hd__buf_4 _15306_ (.A(_07904_),
    .X(_07951_));
 sky130_fd_sc_hd__or3_1 _15307_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_07906_),
    .X(_07952_));
 sky130_fd_sc_hd__o21ai_1 _15308_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_07906_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_07953_));
 sky130_fd_sc_hd__and2_1 _15309_ (.A(_07952_),
    .B(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__mux2_2 _15310_ (.A0(_07954_),
    .A1(\rbzero.debug_overlay.playerY[-4] ),
    .S(_05374_),
    .X(_07955_));
 sky130_fd_sc_hd__nand2_1 _15311_ (.A(_07951_),
    .B(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__a21oi_1 _15312_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_07925_),
    .B1(_05207_),
    .Y(_07957_));
 sky130_fd_sc_hd__a22o_4 _15313_ (.A1(_07945_),
    .A2(_07950_),
    .B1(_07956_),
    .B2(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__buf_4 _15314_ (.A(_07958_),
    .X(_07959_));
 sky130_fd_sc_hd__mux2_1 _15315_ (.A0(_05360_),
    .A1(_05472_),
    .S(\rbzero.wall_tracer.side ),
    .X(_07960_));
 sky130_fd_sc_hd__nand2_1 _15316_ (.A(\rbzero.wall_tracer.state[3] ),
    .B(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__o21ai_4 _15317_ (.A1(_07933_),
    .A2(_07530_),
    .B1(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__a21o_1 _15318_ (.A1(_07903_),
    .A2(\rbzero.wall_tracer.stepDistY[-6] ),
    .B1(_05195_),
    .X(_07963_));
 sky130_fd_sc_hd__a21oi_4 _15319_ (.A1(_04013_),
    .A2(_07962_),
    .B1(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__nor2_2 _15320_ (.A(_05196_),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_07965_));
 sky130_fd_sc_hd__or2_1 _15321_ (.A(_07964_),
    .B(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__clkbuf_4 _15322_ (.A(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__nor2_1 _15323_ (.A(_07959_),
    .B(_07967_),
    .Y(_07968_));
 sky130_fd_sc_hd__xor2_1 _15324_ (.A(_07944_),
    .B(_07968_),
    .X(_07969_));
 sky130_fd_sc_hd__buf_6 _15325_ (.A(\rbzero.wall_tracer.state[3] ),
    .X(_07970_));
 sky130_fd_sc_hd__inv_2 _15326_ (.A(\rbzero.wall_tracer.side ),
    .Y(_07971_));
 sky130_fd_sc_hd__nor2_1 _15327_ (.A(_07971_),
    .B(_05488_),
    .Y(_07972_));
 sky130_fd_sc_hd__a211o_1 _15328_ (.A1(_07971_),
    .A2(_05340_),
    .B1(_07972_),
    .C1(_05193_),
    .X(_07973_));
 sky130_fd_sc_hd__o21ai_4 _15329_ (.A1(_07970_),
    .A2(_07549_),
    .B1(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__nor2_1 _15330_ (.A(_07925_),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_07975_));
 sky130_fd_sc_hd__a211o_2 _15331_ (.A1(_07925_),
    .A2(_07974_),
    .B1(_07975_),
    .C1(_05207_),
    .X(_07976_));
 sky130_fd_sc_hd__a21boi_4 _15332_ (.A1(_05208_),
    .A2(\rbzero.wall_tracer.stepDistX[-2] ),
    .B1_N(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__or2_1 _15333_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_07903_),
    .X(_07978_));
 sky130_fd_sc_hd__o211a_1 _15334_ (.A1(\rbzero.debug_overlay.playerY[-9] ),
    .A2(_04013_),
    .B1(_05196_),
    .C1(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__a21oi_4 _15335_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_05206_),
    .B1(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__clkbuf_4 _15336_ (.A(_07980_),
    .X(_07981_));
 sky130_fd_sc_hd__xor2_1 _15337_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .X(_07982_));
 sky130_fd_sc_hd__mux2_1 _15338_ (.A0(_07982_),
    .A1(\rbzero.debug_overlay.playerY[-8] ),
    .S(_05373_),
    .X(_07983_));
 sky130_fd_sc_hd__mux2_1 _15339_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_07983_),
    .S(_07903_),
    .X(_07984_));
 sky130_fd_sc_hd__xnor2_1 _15340_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_07985_));
 sky130_fd_sc_hd__nor2_1 _15341_ (.A(_05495_),
    .B(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__a211o_1 _15342_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_05496_),
    .B1(_07986_),
    .C1(_05196_),
    .X(_07987_));
 sky130_fd_sc_hd__o21ai_4 _15343_ (.A1(_05206_),
    .A2(_07984_),
    .B1(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__clkbuf_4 _15344_ (.A(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__buf_4 _15345_ (.A(_05196_),
    .X(_07990_));
 sky130_fd_sc_hd__mux2_1 _15346_ (.A0(_05345_),
    .A1(_05466_),
    .S(_07893_),
    .X(_07991_));
 sky130_fd_sc_hd__mux2_2 _15347_ (.A0(_07545_),
    .A1(_07991_),
    .S(\rbzero.wall_tracer.state[3] ),
    .X(_07992_));
 sky130_fd_sc_hd__a21o_1 _15348_ (.A1(_07904_),
    .A2(\rbzero.wall_tracer.stepDistY[-3] ),
    .B1(_05206_),
    .X(_07993_));
 sky130_fd_sc_hd__a21oi_4 _15349_ (.A1(_07925_),
    .A2(_07992_),
    .B1(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__o21bai_4 _15350_ (.A1(_07990_),
    .A2(\rbzero.wall_tracer.stepDistX[-3] ),
    .B1_N(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__clkbuf_4 _15351_ (.A(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__o22ai_1 _15352_ (.A1(_07977_),
    .A2(_07981_),
    .B1(_07989_),
    .B2(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__o21ai_1 _15353_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_07998_));
 sky130_fd_sc_hd__nand2_1 _15354_ (.A(_07897_),
    .B(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__inv_2 _15355_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_08000_));
 sky130_fd_sc_hd__mux2_2 _15356_ (.A0(_07999_),
    .A1(_08000_),
    .S(_05496_),
    .X(_08001_));
 sky130_fd_sc_hd__clkbuf_4 _15357_ (.A(_07904_),
    .X(_08002_));
 sky130_fd_sc_hd__o21ai_1 _15358_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_08003_));
 sky130_fd_sc_hd__and2_1 _15359_ (.A(_07905_),
    .B(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__mux2_2 _15360_ (.A0(_08004_),
    .A1(\rbzero.debug_overlay.playerY[-7] ),
    .S(_05374_),
    .X(_08005_));
 sky130_fd_sc_hd__nand2_1 _15361_ (.A(_08002_),
    .B(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__a21oi_1 _15362_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_04014_),
    .B1(_05207_),
    .Y(_08007_));
 sky130_fd_sc_hd__a22o_4 _15363_ (.A1(_07945_),
    .A2(_08001_),
    .B1(_08006_),
    .B2(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__nor2_1 _15364_ (.A(_08008_),
    .B(_07932_),
    .Y(_08009_));
 sky130_fd_sc_hd__or4_1 _15365_ (.A(_07977_),
    .B(_07995_),
    .C(_07981_),
    .D(_07989_),
    .X(_08010_));
 sky130_fd_sc_hd__a21bo_1 _15366_ (.A1(_07997_),
    .A2(_08009_),
    .B1_N(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__or2b_1 _15367_ (.A(_07969_),
    .B_N(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__xor2_1 _15368_ (.A(_08011_),
    .B(_07969_),
    .X(_08013_));
 sky130_fd_sc_hd__o22ai_1 _15369_ (.A1(_07913_),
    .A2(_07941_),
    .B1(_07967_),
    .B2(_07924_),
    .Y(_08014_));
 sky130_fd_sc_hd__mux2_1 _15370_ (.A0(_05351_),
    .A1(_05475_),
    .S(_07893_),
    .X(_08015_));
 sky130_fd_sc_hd__nand2_1 _15371_ (.A(_07933_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__o21ai_1 _15372_ (.A1(_07933_),
    .A2(_07524_),
    .B1(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__a21o_1 _15373_ (.A1(_07903_),
    .A2(\rbzero.wall_tracer.stepDistY[-7] ),
    .B1(_05195_),
    .X(_08018_));
 sky130_fd_sc_hd__a21oi_2 _15374_ (.A1(_04013_),
    .A2(_08017_),
    .B1(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nor2_1 _15375_ (.A(_05197_),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_08020_));
 sky130_fd_sc_hd__or2_1 _15376_ (.A(_08019_),
    .B(_08020_),
    .X(_08021_));
 sky130_fd_sc_hd__clkbuf_4 _15377_ (.A(_08021_),
    .X(_08022_));
 sky130_fd_sc_hd__nor2_1 _15378_ (.A(_07958_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__or4_1 _15379_ (.A(_07913_),
    .B(_07924_),
    .C(_07941_),
    .D(_07967_),
    .X(_08024_));
 sky130_fd_sc_hd__a21bo_1 _15380_ (.A1(_08014_),
    .A2(_08023_),
    .B1_N(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__or2b_1 _15381_ (.A(_08013_),
    .B_N(_08025_),
    .X(_08026_));
 sky130_fd_sc_hd__or2_1 _15382_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_07946_),
    .X(_08027_));
 sky130_fd_sc_hd__or3_4 _15383_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__or2_1 _15384_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_07952_),
    .X(_08029_));
 sky130_fd_sc_hd__or3_1 _15385_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_08029_),
    .X(_08030_));
 sky130_fd_sc_hd__nor2_1 _15386_ (.A(_05374_),
    .B(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__mux2_1 _15387_ (.A0(\rbzero.wall_tracer.visualWallDist[0] ),
    .A1(_08031_),
    .S(_07904_),
    .X(_08032_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_07990_),
    .B(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__o31a_4 _15389_ (.A1(_07990_),
    .A2(_05496_),
    .A3(_08028_),
    .B1(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__clkbuf_4 _15390_ (.A(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__mux2_1 _15391_ (.A0(_05355_),
    .A1(_05477_),
    .S(_07893_),
    .X(_08036_));
 sky130_fd_sc_hd__mux2_4 _15392_ (.A0(_07502_),
    .A1(_08036_),
    .S(_07933_),
    .X(_08037_));
 sky130_fd_sc_hd__a21o_1 _15393_ (.A1(_07904_),
    .A2(\rbzero.wall_tracer.stepDistY[-9] ),
    .B1(_05206_),
    .X(_08038_));
 sky130_fd_sc_hd__a21o_2 _15394_ (.A1(_07925_),
    .A2(_08037_),
    .B1(_08038_),
    .X(_08039_));
 sky130_fd_sc_hd__or2_1 _15395_ (.A(_05197_),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_08040_));
 sky130_fd_sc_hd__nand2_1 _15396_ (.A(_08039_),
    .B(_08040_),
    .Y(_08041_));
 sky130_fd_sc_hd__clkbuf_4 _15397_ (.A(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__or2_1 _15398_ (.A(_08035_),
    .B(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__nand2_4 _15399_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_07925_),
    .Y(_08044_));
 sky130_fd_sc_hd__or2_1 _15400_ (.A(_07945_),
    .B(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__clkbuf_4 _15401_ (.A(_08045_),
    .X(_08046_));
 sky130_fd_sc_hd__buf_4 _15402_ (.A(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__a211oi_1 _15403_ (.A1(_07486_),
    .A2(_07455_),
    .B1(_07483_),
    .C1(\rbzero.wall_tracer.state[3] ),
    .Y(_08048_));
 sky130_fd_sc_hd__inv_2 _15404_ (.A(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_08049_));
 sky130_fd_sc_hd__nand2_1 _15405_ (.A(\rbzero.wall_tracer.side ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_08050_));
 sky130_fd_sc_hd__o211a_1 _15406_ (.A1(\rbzero.wall_tracer.side ),
    .A2(_08049_),
    .B1(_08050_),
    .C1(\rbzero.wall_tracer.state[3] ),
    .X(_08051_));
 sky130_fd_sc_hd__nand2_1 _15407_ (.A(_07903_),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_08052_));
 sky130_fd_sc_hd__o311a_4 _15408_ (.A1(_07903_),
    .A2(_08048_),
    .A3(_08051_),
    .B1(_08052_),
    .C1(_05196_),
    .X(_08053_));
 sky130_fd_sc_hd__buf_4 _15409_ (.A(_08053_),
    .X(_08054_));
 sky130_fd_sc_hd__nor2_1 _15410_ (.A(_08047_),
    .B(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__xnor2_1 _15411_ (.A(_08043_),
    .B(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__nand2_2 _15412_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_04015_),
    .Y(_08057_));
 sky130_fd_sc_hd__or2_2 _15413_ (.A(_05209_),
    .B(_08057_),
    .X(_08058_));
 sky130_fd_sc_hd__clkbuf_4 _15414_ (.A(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__mux2_1 _15415_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(\rbzero.wall_tracer.side ),
    .X(_08060_));
 sky130_fd_sc_hd__a21o_1 _15416_ (.A1(_07933_),
    .A2(_08060_),
    .B1(_07903_),
    .X(_08061_));
 sky130_fd_sc_hd__a21oi_4 _15417_ (.A1(_05193_),
    .A2(_07465_),
    .B1(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__nor2_1 _15418_ (.A(_08059_),
    .B(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__xor2_1 _15419_ (.A(_08056_),
    .B(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__nand2_1 _15420_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_07946_),
    .Y(_08065_));
 sky130_fd_sc_hd__nand2_1 _15421_ (.A(_08027_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__inv_2 _15422_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_08067_));
 sky130_fd_sc_hd__mux2_1 _15423_ (.A0(_08066_),
    .A1(_08067_),
    .S(_05495_),
    .X(_08068_));
 sky130_fd_sc_hd__nand2_1 _15424_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_07952_),
    .Y(_08069_));
 sky130_fd_sc_hd__and2_1 _15425_ (.A(_08029_),
    .B(_08069_),
    .X(_08070_));
 sky130_fd_sc_hd__mux2_1 _15426_ (.A0(_08070_),
    .A1(\rbzero.debug_overlay.playerY[-3] ),
    .S(_05373_),
    .X(_08071_));
 sky130_fd_sc_hd__nand2_1 _15427_ (.A(_07904_),
    .B(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21oi_1 _15428_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_04013_),
    .B1(_05206_),
    .Y(_08073_));
 sky130_fd_sc_hd__a22o_2 _15429_ (.A1(_05206_),
    .A2(_08068_),
    .B1(_08072_),
    .B2(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__clkbuf_4 _15430_ (.A(_07964_),
    .X(_08075_));
 sky130_fd_sc_hd__or3_1 _15431_ (.A(_08074_),
    .B(_08075_),
    .C(_07965_),
    .X(_08076_));
 sky130_fd_sc_hd__xnor2_1 _15432_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_08027_),
    .Y(_08077_));
 sky130_fd_sc_hd__inv_2 _15433_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .Y(_08078_));
 sky130_fd_sc_hd__mux2_1 _15434_ (.A0(_08077_),
    .A1(_08078_),
    .S(_05496_),
    .X(_08079_));
 sky130_fd_sc_hd__xor2_1 _15435_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_08029_),
    .X(_08080_));
 sky130_fd_sc_hd__mux2_2 _15436_ (.A0(_08080_),
    .A1(\rbzero.debug_overlay.playerY[-2] ),
    .S(_05373_),
    .X(_08081_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(_07951_),
    .B(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__a21oi_1 _15438_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_07925_),
    .B1(_05206_),
    .Y(_08083_));
 sky130_fd_sc_hd__a22o_4 _15439_ (.A1(_05207_),
    .A2(_08079_),
    .B1(_08082_),
    .B2(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__or3_2 _15440_ (.A(_08084_),
    .B(_08019_),
    .C(_08020_),
    .X(_08085_));
 sky130_fd_sc_hd__or2_1 _15441_ (.A(_08076_),
    .B(_08085_),
    .X(_08086_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(_08076_),
    .B(_08085_),
    .Y(_08087_));
 sky130_fd_sc_hd__o21ai_1 _15443_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_08029_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_08088_));
 sky130_fd_sc_hd__and2_1 _15444_ (.A(_08030_),
    .B(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__mux2_2 _15445_ (.A0(_08089_),
    .A1(\rbzero.debug_overlay.playerY[-1] ),
    .S(_05373_),
    .X(_08090_));
 sky130_fd_sc_hd__mux2_1 _15446_ (.A0(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A1(_08090_),
    .S(_07951_),
    .X(_08091_));
 sky130_fd_sc_hd__o21ai_1 _15447_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_08027_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_08092_));
 sky130_fd_sc_hd__and2_1 _15448_ (.A(_08028_),
    .B(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__mux2_1 _15449_ (.A0(_08093_),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_05496_),
    .X(_08094_));
 sky130_fd_sc_hd__or2_1 _15450_ (.A(_05197_),
    .B(_08094_),
    .X(_08095_));
 sky130_fd_sc_hd__o21ai_4 _15451_ (.A1(_07945_),
    .A2(_08091_),
    .B1(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__clkbuf_4 _15452_ (.A(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__o21a_1 _15453_ (.A1(_07893_),
    .A2(_05353_),
    .B1(\rbzero.wall_tracer.state[3] ),
    .X(_08098_));
 sky130_fd_sc_hd__o21ai_2 _15454_ (.A1(_07971_),
    .A2(_05481_),
    .B1(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__o21ai_2 _15455_ (.A1(_07933_),
    .A2(_07514_),
    .B1(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__a21o_1 _15456_ (.A1(_07904_),
    .A2(\rbzero.wall_tracer.stepDistY[-8] ),
    .B1(_05195_),
    .X(_08101_));
 sky130_fd_sc_hd__a21oi_4 _15457_ (.A1(_07925_),
    .A2(_08100_),
    .B1(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__nor2_2 _15458_ (.A(_05197_),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_08103_));
 sky130_fd_sc_hd__or2_4 _15459_ (.A(_08102_),
    .B(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__nor2_1 _15460_ (.A(_08097_),
    .B(_08104_),
    .Y(_08105_));
 sky130_fd_sc_hd__and3_1 _15461_ (.A(_08086_),
    .B(_08087_),
    .C(_08105_),
    .X(_08106_));
 sky130_fd_sc_hd__a21oi_1 _15462_ (.A1(_08086_),
    .A2(_08087_),
    .B1(_08105_),
    .Y(_08107_));
 sky130_fd_sc_hd__or2_1 _15463_ (.A(_08106_),
    .B(_08107_),
    .X(_08108_));
 sky130_fd_sc_hd__clkbuf_4 _15464_ (.A(_08074_),
    .X(_08109_));
 sky130_fd_sc_hd__or3_1 _15465_ (.A(_08109_),
    .B(_08085_),
    .C(_08104_),
    .X(_08110_));
 sky130_fd_sc_hd__buf_4 _15466_ (.A(_08109_),
    .X(_08111_));
 sky130_fd_sc_hd__clkbuf_4 _15467_ (.A(_08102_),
    .X(_08112_));
 sky130_fd_sc_hd__or3_1 _15468_ (.A(_08084_),
    .B(_08112_),
    .C(_08103_),
    .X(_08113_));
 sky130_fd_sc_hd__o21ai_1 _15469_ (.A1(_08111_),
    .A2(_08022_),
    .B1(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_1 _15470_ (.A(_08110_),
    .B(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__or2_1 _15471_ (.A(_08097_),
    .B(_08042_),
    .X(_08116_));
 sky130_fd_sc_hd__o21a_1 _15472_ (.A1(_08115_),
    .A2(_08116_),
    .B1(_08110_),
    .X(_08117_));
 sky130_fd_sc_hd__xor2_1 _15473_ (.A(_08108_),
    .B(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__xnor2_1 _15474_ (.A(_08064_),
    .B(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__a21o_1 _15475_ (.A1(_08012_),
    .A2(_08026_),
    .B1(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__nand3_1 _15476_ (.A(_08012_),
    .B(_08026_),
    .C(_08119_),
    .Y(_08121_));
 sky130_fd_sc_hd__nand2_1 _15477_ (.A(_08120_),
    .B(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__inv_2 _15478_ (.A(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_08123_));
 sky130_fd_sc_hd__a211o_4 _15479_ (.A1(_07951_),
    .A2(_08123_),
    .B1(_08062_),
    .C1(_05207_),
    .X(_08124_));
 sky130_fd_sc_hd__o21bai_4 _15480_ (.A1(_05196_),
    .A2(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1_N(_08053_),
    .Y(_08125_));
 sky130_fd_sc_hd__or4_1 _15481_ (.A(_08034_),
    .B(_08046_),
    .C(_08124_),
    .D(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__inv_2 _15482_ (.A(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__clkbuf_4 _15483_ (.A(_08125_),
    .X(_08128_));
 sky130_fd_sc_hd__clkbuf_4 _15484_ (.A(_08035_),
    .X(_08129_));
 sky130_fd_sc_hd__o22a_1 _15485_ (.A1(_08047_),
    .A2(_08124_),
    .B1(_08128_),
    .B2(_08129_),
    .X(_08130_));
 sky130_fd_sc_hd__nor2_1 _15486_ (.A(_08127_),
    .B(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__mux2_1 _15487_ (.A0(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .S(_07893_),
    .X(_08132_));
 sky130_fd_sc_hd__mux2_1 _15488_ (.A0(_07460_),
    .A1(_08132_),
    .S(_07933_),
    .X(_08133_));
 sky130_fd_sc_hd__or2_1 _15489_ (.A(_04013_),
    .B(\rbzero.wall_tracer.stepDistY[-12] ),
    .X(_08134_));
 sky130_fd_sc_hd__o211ai_4 _15490_ (.A1(_07951_),
    .A2(_08133_),
    .B1(_08134_),
    .C1(_05197_),
    .Y(_08135_));
 sky130_fd_sc_hd__nor2_1 _15491_ (.A(_08059_),
    .B(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__xor2_2 _15492_ (.A(_08131_),
    .B(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__xnor2_1 _15493_ (.A(_08115_),
    .B(_08116_),
    .Y(_08138_));
 sky130_fd_sc_hd__or2_1 _15494_ (.A(_08109_),
    .B(_08042_),
    .X(_08139_));
 sky130_fd_sc_hd__o22a_1 _15495_ (.A1(_08109_),
    .A2(_08104_),
    .B1(_08042_),
    .B2(_08084_),
    .X(_08140_));
 sky130_fd_sc_hd__or2_1 _15496_ (.A(_08097_),
    .B(_08128_),
    .X(_08141_));
 sky130_fd_sc_hd__o22a_1 _15497_ (.A1(_08113_),
    .A2(_08139_),
    .B1(_08140_),
    .B2(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__xor2_1 _15498_ (.A(_08138_),
    .B(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__nor2_1 _15499_ (.A(_08138_),
    .B(_08142_),
    .Y(_08144_));
 sky130_fd_sc_hd__a21o_1 _15500_ (.A1(_08137_),
    .A2(_08143_),
    .B1(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__or2b_1 _15501_ (.A(_08122_),
    .B_N(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__buf_4 _15502_ (.A(_07945_),
    .X(_08147_));
 sky130_fd_sc_hd__buf_6 _15503_ (.A(_04014_),
    .X(_08148_));
 sky130_fd_sc_hd__nand2_4 _15504_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__or2_2 _15505_ (.A(_08147_),
    .B(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__clkbuf_4 _15506_ (.A(_08150_),
    .X(_08151_));
 sky130_fd_sc_hd__or2_1 _15507_ (.A(_08135_),
    .B(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__a21oi_1 _15508_ (.A1(_08131_),
    .A2(_08136_),
    .B1(_08127_),
    .Y(_08153_));
 sky130_fd_sc_hd__or2_1 _15509_ (.A(_08152_),
    .B(_08153_),
    .X(_08154_));
 sky130_fd_sc_hd__and2b_1 _15510_ (.A_N(_08043_),
    .B(_08055_),
    .X(_08155_));
 sky130_fd_sc_hd__and2_1 _15511_ (.A(_08056_),
    .B(_08063_),
    .X(_08156_));
 sky130_fd_sc_hd__nand2_4 _15512_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08148_),
    .Y(_08157_));
 sky130_fd_sc_hd__or2_1 _15513_ (.A(_05208_),
    .B(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__clkbuf_4 _15514_ (.A(_08158_),
    .X(_08159_));
 sky130_fd_sc_hd__clkbuf_4 _15515_ (.A(_08124_),
    .X(_08160_));
 sky130_fd_sc_hd__nor3_1 _15516_ (.A(_08159_),
    .B(_08160_),
    .C(_08152_),
    .Y(_08161_));
 sky130_fd_sc_hd__clkbuf_4 _15517_ (.A(_08135_),
    .X(_08162_));
 sky130_fd_sc_hd__o22a_1 _15518_ (.A1(_08162_),
    .A2(_08159_),
    .B1(_08160_),
    .B2(_08151_),
    .X(_08163_));
 sky130_fd_sc_hd__nor2_1 _15519_ (.A(_08161_),
    .B(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__o21a_1 _15520_ (.A1(_08155_),
    .A2(_08156_),
    .B1(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__nor3_1 _15521_ (.A(_08155_),
    .B(_08156_),
    .C(_08164_),
    .Y(_08166_));
 sky130_fd_sc_hd__nor2_1 _15522_ (.A(_08165_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__xor2_1 _15523_ (.A(_08154_),
    .B(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__a21oi_2 _15524_ (.A1(_08120_),
    .A2(_08146_),
    .B1(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__buf_4 _15525_ (.A(_07981_),
    .X(_08170_));
 sky130_fd_sc_hd__a21oi_4 _15526_ (.A1(_07549_),
    .A2(_07552_),
    .B1(_07555_),
    .Y(_08171_));
 sky130_fd_sc_hd__xnor2_1 _15527_ (.A(_07560_),
    .B(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _15528_ (.A(_07894_),
    .B(_05490_),
    .Y(_08173_));
 sky130_fd_sc_hd__o211a_1 _15529_ (.A1(_07894_),
    .A2(_05342_),
    .B1(_08173_),
    .C1(_07970_),
    .X(_08174_));
 sky130_fd_sc_hd__a211o_1 _15530_ (.A1(_05194_),
    .A2(_08172_),
    .B1(_08174_),
    .C1(_08002_),
    .X(_08175_));
 sky130_fd_sc_hd__o21a_1 _15531_ (.A1(_08148_),
    .A2(\rbzero.wall_tracer.stepDistY[1] ),
    .B1(_07990_),
    .X(_08176_));
 sky130_fd_sc_hd__a22oi_4 _15532_ (.A1(_08147_),
    .A2(\rbzero.wall_tracer.stepDistX[1] ),
    .B1(_08175_),
    .B2(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__clkbuf_4 _15533_ (.A(_08177_),
    .X(_08178_));
 sky130_fd_sc_hd__nor2_1 _15534_ (.A(_08170_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__buf_4 _15535_ (.A(_07989_),
    .X(_08180_));
 sky130_fd_sc_hd__or3_1 _15536_ (.A(_07560_),
    .B(_07562_),
    .C(_08171_),
    .X(_08181_));
 sky130_fd_sc_hd__o21ai_1 _15537_ (.A1(_07560_),
    .A2(_08171_),
    .B1(_07562_),
    .Y(_08182_));
 sky130_fd_sc_hd__a21o_1 _15538_ (.A1(_08181_),
    .A2(_08182_),
    .B1(_07970_),
    .X(_08183_));
 sky130_fd_sc_hd__nor2_1 _15539_ (.A(_07894_),
    .B(_05335_),
    .Y(_08184_));
 sky130_fd_sc_hd__a211o_2 _15540_ (.A1(_07894_),
    .A2(_05456_),
    .B1(_08184_),
    .C1(_05193_),
    .X(_08185_));
 sky130_fd_sc_hd__inv_2 _15541_ (.A(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_08186_));
 sky130_fd_sc_hd__a21o_1 _15542_ (.A1(_07951_),
    .A2(_08186_),
    .B1(_05207_),
    .X(_08187_));
 sky130_fd_sc_hd__a31o_4 _15543_ (.A1(_08148_),
    .A2(_08183_),
    .A3(_08185_),
    .B1(_08187_),
    .X(_08188_));
 sky130_fd_sc_hd__a21boi_4 _15544_ (.A1(_08147_),
    .A2(\rbzero.wall_tracer.stepDistX[2] ),
    .B1_N(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__nor2_1 _15545_ (.A(_08180_),
    .B(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__nor2_1 _15546_ (.A(_08177_),
    .B(_07989_),
    .Y(_08191_));
 sky130_fd_sc_hd__o21ba_1 _15547_ (.A1(_08170_),
    .A2(_08189_),
    .B1_N(_08191_),
    .X(_08192_));
 sky130_fd_sc_hd__a21o_1 _15548_ (.A1(_08179_),
    .A2(_08190_),
    .B1(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__buf_4 _15549_ (.A(_08008_),
    .X(_08194_));
 sky130_fd_sc_hd__nor2_1 _15550_ (.A(_07893_),
    .B(_05369_),
    .Y(_08195_));
 sky130_fd_sc_hd__a211o_1 _15551_ (.A1(_07894_),
    .A2(_05459_),
    .B1(_08195_),
    .C1(_05193_),
    .X(_08196_));
 sky130_fd_sc_hd__and3_1 _15552_ (.A(_07549_),
    .B(_07552_),
    .C(_07555_),
    .X(_08197_));
 sky130_fd_sc_hd__o21ai_1 _15553_ (.A1(_08171_),
    .A2(_08197_),
    .B1(_05193_),
    .Y(_08198_));
 sky130_fd_sc_hd__a21o_2 _15554_ (.A1(_08196_),
    .A2(_08198_),
    .B1(_07951_),
    .X(_08199_));
 sky130_fd_sc_hd__inv_2 _15555_ (.A(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_08200_));
 sky130_fd_sc_hd__a21oi_2 _15556_ (.A1(_08002_),
    .A2(_08200_),
    .B1(_07945_),
    .Y(_08201_));
 sky130_fd_sc_hd__nand2_4 _15557_ (.A(_08199_),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_2 _15558_ (.A(_05208_),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_08203_));
 sky130_fd_sc_hd__and2_2 _15559_ (.A(_08202_),
    .B(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__nor2_2 _15560_ (.A(_08194_),
    .B(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__xnor2_4 _15561_ (.A(_08193_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__inv_2 _15562_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_08207_));
 sky130_fd_sc_hd__nor4_2 _15563_ (.A(_07560_),
    .B(_07562_),
    .C(_07564_),
    .D(_08171_),
    .Y(_08208_));
 sky130_fd_sc_hd__o31a_1 _15564_ (.A1(_07560_),
    .A2(_07562_),
    .A3(_08171_),
    .B1(_07564_),
    .X(_08209_));
 sky130_fd_sc_hd__o21ai_1 _15565_ (.A1(_08208_),
    .A2(_08209_),
    .B1(_05194_),
    .Y(_08210_));
 sky130_fd_sc_hd__nand2_1 _15566_ (.A(_07894_),
    .B(_05454_),
    .Y(_08211_));
 sky130_fd_sc_hd__o211a_1 _15567_ (.A1(_07894_),
    .A2(_05331_),
    .B1(_08211_),
    .C1(_07970_),
    .X(_08212_));
 sky130_fd_sc_hd__nor2_1 _15568_ (.A(_08002_),
    .B(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__a221o_1 _15569_ (.A1(_08002_),
    .A2(_08207_),
    .B1(_08210_),
    .B2(_08213_),
    .C1(_07945_),
    .X(_08214_));
 sky130_fd_sc_hd__nand2_8 _15570_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_04012_),
    .Y(_08215_));
 sky130_fd_sc_hd__nor2_2 _15571_ (.A(_08214_),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__and2_1 _15572_ (.A(_08002_),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_08217_));
 sky130_fd_sc_hd__inv_2 _15573_ (.A(_07566_),
    .Y(_08218_));
 sky130_fd_sc_hd__nand2_1 _15574_ (.A(_08218_),
    .B(_08208_),
    .Y(_08219_));
 sky130_fd_sc_hd__or4_1 _15575_ (.A(_07560_),
    .B(_07562_),
    .C(_07564_),
    .D(_08171_),
    .X(_08220_));
 sky130_fd_sc_hd__a21oi_1 _15576_ (.A1(_07566_),
    .A2(_08220_),
    .B1(_07970_),
    .Y(_08221_));
 sky130_fd_sc_hd__nand2_1 _15577_ (.A(_07894_),
    .B(_05494_),
    .Y(_08222_));
 sky130_fd_sc_hd__or2_2 _15578_ (.A(_07893_),
    .B(_05372_),
    .X(_08223_));
 sky130_fd_sc_hd__a31o_2 _15579_ (.A1(_07970_),
    .A2(_08222_),
    .A3(_08223_),
    .B1(_07951_),
    .X(_08224_));
 sky130_fd_sc_hd__a21oi_2 _15580_ (.A1(_08219_),
    .A2(_08221_),
    .B1(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__nand2_4 _15581_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_04012_),
    .Y(_08226_));
 sky130_fd_sc_hd__nor2_4 _15582_ (.A(_05207_),
    .B(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__o21a_1 _15583_ (.A1(_08217_),
    .A2(_08225_),
    .B1(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__xnor2_4 _15584_ (.A(_08216_),
    .B(_08228_),
    .Y(_08229_));
 sky130_fd_sc_hd__clkbuf_4 _15585_ (.A(_08002_),
    .X(_08230_));
 sky130_fd_sc_hd__nand2_1 _15586_ (.A(_08230_),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_08231_));
 sky130_fd_sc_hd__inv_2 _15587_ (.A(_07568_),
    .Y(_08232_));
 sky130_fd_sc_hd__a21oi_1 _15588_ (.A1(_08218_),
    .A2(_08208_),
    .B1(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__and3_1 _15589_ (.A(_08218_),
    .B(_08232_),
    .C(_08208_),
    .X(_08234_));
 sky130_fd_sc_hd__a31oi_4 _15590_ (.A1(_07970_),
    .A2(_08222_),
    .A3(_08223_),
    .B1(_08002_),
    .Y(_08235_));
 sky130_fd_sc_hd__o31ai_2 _15591_ (.A1(_07970_),
    .A2(_08233_),
    .A3(_08234_),
    .B1(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__a21o_2 _15592_ (.A1(_08231_),
    .A2(_08236_),
    .B1(_05209_),
    .X(_08237_));
 sky130_fd_sc_hd__nand2_4 _15593_ (.A(\rbzero.wall_tracer.visualWallDist[-12] ),
    .B(_04014_),
    .Y(_08238_));
 sky130_fd_sc_hd__clkbuf_4 _15594_ (.A(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__nor2_2 _15595_ (.A(_08237_),
    .B(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__xor2_4 _15596_ (.A(_08229_),
    .B(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__o21ai_4 _15597_ (.A1(_08217_),
    .A2(_08225_),
    .B1(_05198_),
    .Y(_08242_));
 sky130_fd_sc_hd__a2111o_1 _15598_ (.A1(_08210_),
    .A2(_08213_),
    .B1(_07598_),
    .C1(_08002_),
    .D1(_05208_),
    .X(_08243_));
 sky130_fd_sc_hd__a2111o_1 _15599_ (.A1(_08183_),
    .A2(_08185_),
    .B1(_07602_),
    .C1(_08230_),
    .D1(_05208_),
    .X(_08244_));
 sky130_fd_sc_hd__xnor2_1 _15600_ (.A(_08243_),
    .B(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__or2_1 _15601_ (.A(_08243_),
    .B(_08244_),
    .X(_08246_));
 sky130_fd_sc_hd__o31a_2 _15602_ (.A1(_08242_),
    .A2(_08239_),
    .A3(_08245_),
    .B1(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__xor2_4 _15603_ (.A(_08241_),
    .B(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__xnor2_4 _15604_ (.A(_08206_),
    .B(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__nor2_4 _15605_ (.A(_07945_),
    .B(_08238_),
    .Y(_08250_));
 sky130_fd_sc_hd__o21a_1 _15606_ (.A1(_08217_),
    .A2(_08225_),
    .B1(_08250_),
    .X(_08251_));
 sky130_fd_sc_hd__xor2_1 _15607_ (.A(_08245_),
    .B(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__a2111o_1 _15608_ (.A1(_08183_),
    .A2(_08185_),
    .B1(_07598_),
    .C1(_08002_),
    .D1(_05208_),
    .X(_08253_));
 sky130_fd_sc_hd__a21o_1 _15609_ (.A1(_05193_),
    .A2(_08172_),
    .B1(_08174_),
    .X(_08254_));
 sky130_fd_sc_hd__and4_1 _15610_ (.A(_07601_),
    .B(_04015_),
    .C(_05198_),
    .D(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__xnor2_1 _15611_ (.A(_08253_),
    .B(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__clkbuf_4 _15612_ (.A(_08214_),
    .X(_08257_));
 sky130_fd_sc_hd__nor2_1 _15613_ (.A(_08257_),
    .B(_08238_),
    .Y(_08258_));
 sky130_fd_sc_hd__nand2_4 _15614_ (.A(_08175_),
    .B(_08176_),
    .Y(_08259_));
 sky130_fd_sc_hd__or3_1 _15615_ (.A(_08259_),
    .B(_08226_),
    .C(_08244_),
    .X(_08260_));
 sky130_fd_sc_hd__a21boi_1 _15616_ (.A1(_08256_),
    .A2(_08258_),
    .B1_N(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__xor2_1 _15617_ (.A(_08252_),
    .B(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__a21o_2 _15618_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_08147_),
    .B1(_07979_),
    .X(_08263_));
 sky130_fd_sc_hd__a21bo_2 _15619_ (.A1(_08199_),
    .A2(_08201_),
    .B1_N(_08203_),
    .X(_08264_));
 sky130_fd_sc_hd__and2_1 _15620_ (.A(_08263_),
    .B(_08264_),
    .X(_08265_));
 sky130_fd_sc_hd__clkinv_2 _15621_ (.A(_07988_),
    .Y(_08266_));
 sky130_fd_sc_hd__a2bb2o_1 _15622_ (.A1_N(_07981_),
    .A2_N(_08177_),
    .B1(_08266_),
    .B2(_08264_),
    .X(_08267_));
 sky130_fd_sc_hd__a21bo_1 _15623_ (.A1(_08191_),
    .A2(_08265_),
    .B1_N(_08267_),
    .X(_08268_));
 sky130_fd_sc_hd__inv_2 _15624_ (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_08269_));
 sky130_fd_sc_hd__inv_2 _15625_ (.A(_07551_),
    .Y(_08270_));
 sky130_fd_sc_hd__a22o_1 _15626_ (.A1(_07487_),
    .A2(_07455_),
    .B1(_07548_),
    .B2(_07551_),
    .X(_08271_));
 sky130_fd_sc_hd__a211o_2 _15627_ (.A1(_07549_),
    .A2(_08270_),
    .B1(_08271_),
    .C1(_07933_),
    .X(_08272_));
 sky130_fd_sc_hd__mux2_1 _15628_ (.A0(_05364_),
    .A1(_05461_),
    .S(_07893_),
    .X(_08273_));
 sky130_fd_sc_hd__o21a_1 _15629_ (.A1(_05193_),
    .A2(_08273_),
    .B1(_04013_),
    .X(_08274_));
 sky130_fd_sc_hd__a22oi_4 _15630_ (.A1(_07951_),
    .A2(\rbzero.wall_tracer.stepDistY[-1] ),
    .B1(_08272_),
    .B2(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__mux2_2 _15631_ (.A0(_08269_),
    .A1(_08275_),
    .S(_07990_),
    .X(_08276_));
 sky130_fd_sc_hd__nor2_1 _15632_ (.A(_08276_),
    .B(_08008_),
    .Y(_08277_));
 sky130_fd_sc_hd__xnor2_1 _15633_ (.A(_08268_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__nor2_1 _15634_ (.A(_08252_),
    .B(_08261_),
    .Y(_08279_));
 sky130_fd_sc_hd__a21oi_2 _15635_ (.A1(_08262_),
    .A2(_08278_),
    .B1(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__xor2_4 _15636_ (.A(_08249_),
    .B(_08280_),
    .X(_08281_));
 sky130_fd_sc_hd__clkbuf_4 _15637_ (.A(_07977_),
    .X(_08282_));
 sky130_fd_sc_hd__buf_4 _15638_ (.A(_07913_),
    .X(_08283_));
 sky130_fd_sc_hd__buf_6 _15639_ (.A(_07924_),
    .X(_08284_));
 sky130_fd_sc_hd__o22ai_1 _15640_ (.A1(_08282_),
    .A2(_08283_),
    .B1(_08284_),
    .B2(_07996_),
    .Y(_08285_));
 sky130_fd_sc_hd__nor2_1 _15641_ (.A(_07959_),
    .B(_07932_),
    .Y(_08286_));
 sky130_fd_sc_hd__or4_1 _15642_ (.A(_07977_),
    .B(_07913_),
    .C(_07924_),
    .D(_07995_),
    .X(_08287_));
 sky130_fd_sc_hd__a21bo_1 _15643_ (.A1(_08285_),
    .A2(_08286_),
    .B1_N(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__a22o_1 _15644_ (.A1(_08191_),
    .A2(_08265_),
    .B1(_08277_),
    .B2(_08267_),
    .X(_08289_));
 sky130_fd_sc_hd__nor2_1 _15645_ (.A(_07977_),
    .B(_07923_),
    .Y(_08290_));
 sky130_fd_sc_hd__nor2_1 _15646_ (.A(_07912_),
    .B(_08276_),
    .Y(_08291_));
 sky130_fd_sc_hd__xnor2_1 _15647_ (.A(_08290_),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__nor2_1 _15648_ (.A(_07996_),
    .B(_07958_),
    .Y(_08293_));
 sky130_fd_sc_hd__xnor2_2 _15649_ (.A(_08292_),
    .B(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__xnor2_2 _15650_ (.A(_08289_),
    .B(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__xnor2_4 _15651_ (.A(_08288_),
    .B(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__xnor2_4 _15652_ (.A(_08281_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__xnor2_1 _15653_ (.A(_08262_),
    .B(_08278_),
    .Y(_08298_));
 sky130_fd_sc_hd__xnor2_1 _15654_ (.A(_08256_),
    .B(_08258_),
    .Y(_08299_));
 sky130_fd_sc_hd__and4_1 _15655_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08148_),
    .C(_05198_),
    .D(_08254_),
    .X(_08300_));
 sky130_fd_sc_hd__and4_1 _15656_ (.A(_07601_),
    .B(_08148_),
    .C(_05198_),
    .D(_08199_),
    .X(_08301_));
 sky130_fd_sc_hd__xnor2_1 _15657_ (.A(_08300_),
    .B(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__and4_1 _15658_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08148_),
    .C(_05198_),
    .D(_08199_),
    .X(_08303_));
 sky130_fd_sc_hd__nand2_1 _15659_ (.A(_08255_),
    .B(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__o31a_1 _15660_ (.A1(_08188_),
    .A2(_08239_),
    .A3(_08302_),
    .B1(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__xor2_1 _15661_ (.A(_08299_),
    .B(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__nor2_1 _15662_ (.A(_08276_),
    .B(_07989_),
    .Y(_08307_));
 sky130_fd_sc_hd__xnor2_1 _15663_ (.A(_08265_),
    .B(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(_08282_),
    .B(_08194_),
    .Y(_08309_));
 sky130_fd_sc_hd__xnor2_2 _15665_ (.A(_08308_),
    .B(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__nor2_1 _15666_ (.A(_08299_),
    .B(_08305_),
    .Y(_08311_));
 sky130_fd_sc_hd__a21oi_1 _15667_ (.A1(_08306_),
    .A2(_08310_),
    .B1(_08311_),
    .Y(_08312_));
 sky130_fd_sc_hd__xor2_1 _15668_ (.A(_08298_),
    .B(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__o22ai_1 _15669_ (.A1(_07913_),
    .A2(_07996_),
    .B1(_07932_),
    .B2(_07924_),
    .Y(_08314_));
 sky130_fd_sc_hd__nor2_1 _15670_ (.A(_07959_),
    .B(_07941_),
    .Y(_08315_));
 sky130_fd_sc_hd__or4_1 _15671_ (.A(_07913_),
    .B(_07924_),
    .C(_07995_),
    .D(_07932_),
    .X(_08316_));
 sky130_fd_sc_hd__a21bo_1 _15672_ (.A1(_08314_),
    .A2(_08315_),
    .B1_N(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__a21o_1 _15673_ (.A1(_08263_),
    .A2(_08264_),
    .B1(_08307_),
    .X(_08318_));
 sky130_fd_sc_hd__and3_1 _15674_ (.A(_08263_),
    .B(_08264_),
    .C(_08307_),
    .X(_08319_));
 sky130_fd_sc_hd__a21o_1 _15675_ (.A1(_08318_),
    .A2(_08309_),
    .B1(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__nand2_1 _15676_ (.A(_08287_),
    .B(_08285_),
    .Y(_08321_));
 sky130_fd_sc_hd__xnor2_1 _15677_ (.A(_08321_),
    .B(_08286_),
    .Y(_08322_));
 sky130_fd_sc_hd__xnor2_1 _15678_ (.A(_08320_),
    .B(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__xnor2_1 _15679_ (.A(_08317_),
    .B(_08323_),
    .Y(_08324_));
 sky130_fd_sc_hd__nor2_1 _15680_ (.A(_08298_),
    .B(_08312_),
    .Y(_08325_));
 sky130_fd_sc_hd__a21oi_2 _15681_ (.A1(_08313_),
    .A2(_08324_),
    .B1(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__xor2_4 _15682_ (.A(_08297_),
    .B(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__a21oi_4 _15683_ (.A1(_08148_),
    .A2(_08037_),
    .B1(_08038_),
    .Y(_08328_));
 sky130_fd_sc_hd__buf_4 _15684_ (.A(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__or4_1 _15685_ (.A(_08035_),
    .B(_08046_),
    .C(_08329_),
    .D(_08104_),
    .X(_08330_));
 sky130_fd_sc_hd__buf_4 _15686_ (.A(_08039_),
    .X(_08331_));
 sky130_fd_sc_hd__nor2_2 _15687_ (.A(_05210_),
    .B(_08044_),
    .Y(_08332_));
 sky130_fd_sc_hd__a2bb2o_1 _15688_ (.A1_N(_08129_),
    .A2_N(_08104_),
    .B1(_08331_),
    .B2(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__nand2_1 _15689_ (.A(_08330_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__clkbuf_4 _15690_ (.A(_08054_),
    .X(_08335_));
 sky130_fd_sc_hd__nor2_1 _15691_ (.A(_08059_),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__xnor2_1 _15692_ (.A(_08334_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__or3_1 _15693_ (.A(_07938_),
    .B(_07939_),
    .C(_08109_),
    .X(_08338_));
 sky130_fd_sc_hd__or3_1 _15694_ (.A(_08084_),
    .B(_07964_),
    .C(_07965_),
    .X(_08339_));
 sky130_fd_sc_hd__or2_1 _15695_ (.A(_08338_),
    .B(_08339_),
    .X(_08340_));
 sky130_fd_sc_hd__nand2_1 _15696_ (.A(_08338_),
    .B(_08339_),
    .Y(_08341_));
 sky130_fd_sc_hd__nor2_1 _15697_ (.A(_08097_),
    .B(_08022_),
    .Y(_08342_));
 sky130_fd_sc_hd__and3_1 _15698_ (.A(_08340_),
    .B(_08341_),
    .C(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__a21oi_1 _15699_ (.A1(_08340_),
    .A2(_08341_),
    .B1(_08342_),
    .Y(_08344_));
 sky130_fd_sc_hd__or2_1 _15700_ (.A(_08343_),
    .B(_08344_),
    .X(_08345_));
 sky130_fd_sc_hd__o21ba_1 _15701_ (.A1(_08076_),
    .A2(_08085_),
    .B1_N(_08106_),
    .X(_08346_));
 sky130_fd_sc_hd__xor2_1 _15702_ (.A(_08345_),
    .B(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__nor2_1 _15703_ (.A(_08345_),
    .B(_08346_),
    .Y(_08348_));
 sky130_fd_sc_hd__a21o_1 _15704_ (.A1(_08337_),
    .A2(_08347_),
    .B1(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__nand2_1 _15705_ (.A(_08320_),
    .B(_08322_),
    .Y(_08350_));
 sky130_fd_sc_hd__or2b_1 _15706_ (.A(_08323_),
    .B_N(_08317_),
    .X(_08351_));
 sky130_fd_sc_hd__or4_1 _15707_ (.A(_08022_),
    .B(_08034_),
    .C(_08045_),
    .D(_08112_),
    .X(_08352_));
 sky130_fd_sc_hd__o22ai_1 _15708_ (.A1(_08022_),
    .A2(_08035_),
    .B1(_08046_),
    .B2(_08112_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_1 _15709_ (.A(_08352_),
    .B(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__or3_1 _15710_ (.A(_08354_),
    .B(_08329_),
    .C(_08058_),
    .X(_08355_));
 sky130_fd_sc_hd__buf_4 _15711_ (.A(_08059_),
    .X(_08356_));
 sky130_fd_sc_hd__o21ai_1 _15712_ (.A1(_08329_),
    .A2(_08356_),
    .B1(_08354_),
    .Y(_08357_));
 sky130_fd_sc_hd__and2_1 _15713_ (.A(_08355_),
    .B(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__nor2_1 _15714_ (.A(_07940_),
    .B(_08084_),
    .Y(_08359_));
 sky130_fd_sc_hd__nor2_1 _15715_ (.A(_07931_),
    .B(_08109_),
    .Y(_08360_));
 sky130_fd_sc_hd__xnor2_1 _15716_ (.A(_08359_),
    .B(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__or2_1 _15717_ (.A(_07967_),
    .B(_08097_),
    .X(_08362_));
 sky130_fd_sc_hd__xnor2_1 _15718_ (.A(_08361_),
    .B(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__o21ba_1 _15719_ (.A1(_08338_),
    .A2(_08339_),
    .B1_N(_08343_),
    .X(_08364_));
 sky130_fd_sc_hd__xor2_1 _15720_ (.A(_08363_),
    .B(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__xnor2_1 _15721_ (.A(_08358_),
    .B(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__a21o_1 _15722_ (.A1(_08350_),
    .A2(_08351_),
    .B1(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__nand3_1 _15723_ (.A(_08350_),
    .B(_08351_),
    .C(_08366_),
    .Y(_08368_));
 sky130_fd_sc_hd__nand2_1 _15724_ (.A(_08367_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__xnor2_2 _15725_ (.A(_08349_),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__xnor2_2 _15726_ (.A(_08327_),
    .B(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__xnor2_1 _15727_ (.A(_08313_),
    .B(_08324_),
    .Y(_08372_));
 sky130_fd_sc_hd__xnor2_1 _15728_ (.A(_08306_),
    .B(_08310_),
    .Y(_08373_));
 sky130_fd_sc_hd__nor2_1 _15729_ (.A(_08188_),
    .B(_08238_),
    .Y(_08374_));
 sky130_fd_sc_hd__xor2_1 _15730_ (.A(_08302_),
    .B(_08374_),
    .X(_08375_));
 sky130_fd_sc_hd__or2_1 _15731_ (.A(_05206_),
    .B(_08215_),
    .X(_08376_));
 sky130_fd_sc_hd__buf_4 _15732_ (.A(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__nor2_1 _15733_ (.A(_08275_),
    .B(_08377_),
    .Y(_08378_));
 sky130_fd_sc_hd__xnor2_2 _15734_ (.A(_08303_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand2_1 _15735_ (.A(_08303_),
    .B(_08378_),
    .Y(_08380_));
 sky130_fd_sc_hd__o31a_1 _15736_ (.A1(_08259_),
    .A2(_08238_),
    .A3(_08379_),
    .B1(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__xor2_1 _15737_ (.A(_08375_),
    .B(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__clkbuf_4 _15738_ (.A(_08276_),
    .X(_08383_));
 sky130_fd_sc_hd__o22ai_1 _15739_ (.A1(_08383_),
    .A2(_07981_),
    .B1(_08180_),
    .B2(_08282_),
    .Y(_08384_));
 sky130_fd_sc_hd__or4_1 _15740_ (.A(_07977_),
    .B(_08276_),
    .C(_07981_),
    .D(_07989_),
    .X(_08385_));
 sky130_fd_sc_hd__nand2_1 _15741_ (.A(_08384_),
    .B(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__nor2_1 _15742_ (.A(_07996_),
    .B(_08194_),
    .Y(_08387_));
 sky130_fd_sc_hd__xnor2_1 _15743_ (.A(_08386_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__nor2_1 _15744_ (.A(_08375_),
    .B(_08381_),
    .Y(_08389_));
 sky130_fd_sc_hd__a21o_1 _15745_ (.A1(_08382_),
    .A2(_08388_),
    .B1(_08389_),
    .X(_08390_));
 sky130_fd_sc_hd__xnor2_1 _15746_ (.A(_08373_),
    .B(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__a21bo_1 _15747_ (.A1(_07943_),
    .A2(_07968_),
    .B1_N(_07942_),
    .X(_08392_));
 sky130_fd_sc_hd__o31a_1 _15748_ (.A1(_07996_),
    .A2(_08194_),
    .A3(_08386_),
    .B1(_08385_),
    .X(_08393_));
 sky130_fd_sc_hd__nand2_1 _15749_ (.A(_08316_),
    .B(_08314_),
    .Y(_08394_));
 sky130_fd_sc_hd__xor2_1 _15750_ (.A(_08394_),
    .B(_08315_),
    .X(_08395_));
 sky130_fd_sc_hd__xnor2_1 _15751_ (.A(_08393_),
    .B(_08395_),
    .Y(_08396_));
 sky130_fd_sc_hd__xnor2_2 _15752_ (.A(_08392_),
    .B(_08396_),
    .Y(_08397_));
 sky130_fd_sc_hd__and2b_1 _15753_ (.A_N(_08373_),
    .B(_08390_),
    .X(_08398_));
 sky130_fd_sc_hd__a21oi_2 _15754_ (.A1(_08391_),
    .A2(_08397_),
    .B1(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__xor2_1 _15755_ (.A(_08372_),
    .B(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__nor2_1 _15756_ (.A(_08108_),
    .B(_08117_),
    .Y(_08401_));
 sky130_fd_sc_hd__a21o_1 _15757_ (.A1(_08064_),
    .A2(_08118_),
    .B1(_08401_),
    .X(_08402_));
 sky130_fd_sc_hd__or2_1 _15758_ (.A(_08393_),
    .B(_08395_),
    .X(_08403_));
 sky130_fd_sc_hd__or2b_1 _15759_ (.A(_08396_),
    .B_N(_08392_),
    .X(_08404_));
 sky130_fd_sc_hd__xnor2_1 _15760_ (.A(_08337_),
    .B(_08347_),
    .Y(_08405_));
 sky130_fd_sc_hd__a21o_1 _15761_ (.A1(_08403_),
    .A2(_08404_),
    .B1(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__nand3_1 _15762_ (.A(_08403_),
    .B(_08404_),
    .C(_08405_),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_1 _15763_ (.A(_08406_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__xnor2_1 _15764_ (.A(_08402_),
    .B(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_08372_),
    .B(_08399_),
    .Y(_08410_));
 sky130_fd_sc_hd__a21oi_2 _15766_ (.A1(_08400_),
    .A2(_08409_),
    .B1(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__xor2_2 _15767_ (.A(_08371_),
    .B(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__or2b_1 _15768_ (.A(_08154_),
    .B_N(_08167_),
    .X(_08413_));
 sky130_fd_sc_hd__or2b_1 _15769_ (.A(_08408_),
    .B_N(_08402_),
    .X(_08414_));
 sky130_fd_sc_hd__or3_1 _15770_ (.A(_08059_),
    .B(_08334_),
    .C(_08335_),
    .X(_08415_));
 sky130_fd_sc_hd__inv_2 _15771_ (.A(_08124_),
    .Y(_08416_));
 sky130_fd_sc_hd__nor2_1 _15772_ (.A(_05208_),
    .B(_08157_),
    .Y(_08417_));
 sky130_fd_sc_hd__nor2_2 _15773_ (.A(_05208_),
    .B(_08149_),
    .Y(_08418_));
 sky130_fd_sc_hd__nand2_1 _15774_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__nor2_1 _15775_ (.A(_08054_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__o22a_1 _15776_ (.A1(_08062_),
    .A2(_08158_),
    .B1(_08150_),
    .B2(_08054_),
    .X(_08421_));
 sky130_fd_sc_hd__a21o_1 _15777_ (.A1(_08416_),
    .A2(_08420_),
    .B1(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__nand2_8 _15778_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_04014_),
    .Y(_08423_));
 sky130_fd_sc_hd__or2_1 _15779_ (.A(_05208_),
    .B(_08423_),
    .X(_08424_));
 sky130_fd_sc_hd__clkbuf_2 _15780_ (.A(_08424_),
    .X(_08425_));
 sky130_fd_sc_hd__or3_1 _15781_ (.A(_08135_),
    .B(_08422_),
    .C(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__clkbuf_4 _15782_ (.A(_08425_),
    .X(_08427_));
 sky130_fd_sc_hd__o21ai_1 _15783_ (.A1(_08135_),
    .A2(_08427_),
    .B1(_08422_),
    .Y(_08428_));
 sky130_fd_sc_hd__nand2_1 _15784_ (.A(_08426_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__and3_1 _15785_ (.A(_08330_),
    .B(_08415_),
    .C(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__a21oi_1 _15786_ (.A1(_08330_),
    .A2(_08415_),
    .B1(_08429_),
    .Y(_08431_));
 sky130_fd_sc_hd__nor2_1 _15787_ (.A(_08430_),
    .B(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__or2_1 _15788_ (.A(_08161_),
    .B(_08165_),
    .X(_08433_));
 sky130_fd_sc_hd__xnor2_1 _15789_ (.A(_08432_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__a21o_1 _15790_ (.A1(_08406_),
    .A2(_08414_),
    .B1(_08434_),
    .X(_08435_));
 sky130_fd_sc_hd__nand3_1 _15791_ (.A(_08406_),
    .B(_08414_),
    .C(_08434_),
    .Y(_08436_));
 sky130_fd_sc_hd__and2_1 _15792_ (.A(_08435_),
    .B(_08436_),
    .X(_08437_));
 sky130_fd_sc_hd__xnor2_2 _15793_ (.A(_08413_),
    .B(_08437_),
    .Y(_08438_));
 sky130_fd_sc_hd__xnor2_2 _15794_ (.A(_08412_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__xnor2_1 _15795_ (.A(_08400_),
    .B(_08409_),
    .Y(_08440_));
 sky130_fd_sc_hd__xnor2_1 _15796_ (.A(_08391_),
    .B(_08397_),
    .Y(_08441_));
 sky130_fd_sc_hd__xnor2_1 _15797_ (.A(_08382_),
    .B(_08388_),
    .Y(_08442_));
 sky130_fd_sc_hd__nor2_1 _15798_ (.A(_08259_),
    .B(_08238_),
    .Y(_08443_));
 sky130_fd_sc_hd__xor2_2 _15799_ (.A(_08379_),
    .B(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__a22o_4 _15800_ (.A1(_07904_),
    .A2(\rbzero.wall_tracer.stepDistY[-1] ),
    .B1(_08272_),
    .B2(_08274_),
    .X(_08445_));
 sky130_fd_sc_hd__nand2_1 _15801_ (.A(_08445_),
    .B(_08227_),
    .Y(_08446_));
 sky130_fd_sc_hd__or2_1 _15802_ (.A(_07974_),
    .B(_08376_),
    .X(_08447_));
 sky130_fd_sc_hd__xnor2_2 _15803_ (.A(_08446_),
    .B(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__or3_1 _15804_ (.A(_08202_),
    .B(_08238_),
    .C(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__o31a_1 _15805_ (.A1(_07976_),
    .A2(_08215_),
    .A3(_08446_),
    .B1(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__xor2_2 _15806_ (.A(_08444_),
    .B(_08450_),
    .X(_08451_));
 sky130_fd_sc_hd__nand2_1 _15807_ (.A(_08010_),
    .B(_07997_),
    .Y(_08452_));
 sky130_fd_sc_hd__xnor2_2 _15808_ (.A(_08452_),
    .B(_08009_),
    .Y(_08453_));
 sky130_fd_sc_hd__nor2_1 _15809_ (.A(_08444_),
    .B(_08450_),
    .Y(_08454_));
 sky130_fd_sc_hd__a21oi_1 _15810_ (.A1(_08451_),
    .A2(_08453_),
    .B1(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__xor2_1 _15811_ (.A(_08442_),
    .B(_08455_),
    .X(_08456_));
 sky130_fd_sc_hd__xnor2_1 _15812_ (.A(_08025_),
    .B(_08013_),
    .Y(_08457_));
 sky130_fd_sc_hd__nor2_1 _15813_ (.A(_08442_),
    .B(_08455_),
    .Y(_08458_));
 sky130_fd_sc_hd__a21oi_1 _15814_ (.A1(_08456_),
    .A2(_08457_),
    .B1(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__xor2_1 _15815_ (.A(_08441_),
    .B(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__xnor2_1 _15816_ (.A(_08145_),
    .B(_08122_),
    .Y(_08461_));
 sky130_fd_sc_hd__nor2_1 _15817_ (.A(_08441_),
    .B(_08459_),
    .Y(_08462_));
 sky130_fd_sc_hd__a21oi_1 _15818_ (.A1(_08460_),
    .A2(_08461_),
    .B1(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand2_1 _15819_ (.A(_08440_),
    .B(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__and3_1 _15820_ (.A(_08120_),
    .B(_08146_),
    .C(_08168_),
    .X(_08465_));
 sky130_fd_sc_hd__nor2_2 _15821_ (.A(_08169_),
    .B(_08465_),
    .Y(_08466_));
 sky130_fd_sc_hd__nor2_1 _15822_ (.A(_08440_),
    .B(_08463_),
    .Y(_08467_));
 sky130_fd_sc_hd__a21oi_2 _15823_ (.A1(_08464_),
    .A2(_08466_),
    .B1(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__xor2_2 _15824_ (.A(_08439_),
    .B(_08468_),
    .X(_08469_));
 sky130_fd_sc_hd__xnor2_2 _15825_ (.A(_08169_),
    .B(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__nand2_1 _15826_ (.A(_08024_),
    .B(_08014_),
    .Y(_08471_));
 sky130_fd_sc_hd__xor2_2 _15827_ (.A(_08471_),
    .B(_08023_),
    .X(_08472_));
 sky130_fd_sc_hd__o22ai_2 _15828_ (.A1(_07995_),
    .A2(_07981_),
    .B1(_07989_),
    .B2(_07931_),
    .Y(_08473_));
 sky130_fd_sc_hd__nor2_1 _15829_ (.A(_08008_),
    .B(_07941_),
    .Y(_08474_));
 sky130_fd_sc_hd__or3_2 _15830_ (.A(_07980_),
    .B(_07929_),
    .C(_07930_),
    .X(_08475_));
 sky130_fd_sc_hd__or3_1 _15831_ (.A(_07995_),
    .B(_07989_),
    .C(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__a21bo_1 _15832_ (.A1(_08473_),
    .A2(_08474_),
    .B1_N(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__or2b_1 _15833_ (.A(_08472_),
    .B_N(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__xor2_2 _15834_ (.A(_08477_),
    .B(_08472_),
    .X(_08479_));
 sky130_fd_sc_hd__o22ai_1 _15835_ (.A1(_07913_),
    .A2(_07967_),
    .B1(_08022_),
    .B2(_07923_),
    .Y(_08480_));
 sky130_fd_sc_hd__nor2_1 _15836_ (.A(_07958_),
    .B(_08104_),
    .Y(_08481_));
 sky130_fd_sc_hd__or3_1 _15837_ (.A(_07912_),
    .B(_08019_),
    .C(_08020_),
    .X(_08482_));
 sky130_fd_sc_hd__or3_1 _15838_ (.A(_07923_),
    .B(_07967_),
    .C(_08482_),
    .X(_08483_));
 sky130_fd_sc_hd__a21bo_1 _15839_ (.A1(_08480_),
    .A2(_08481_),
    .B1_N(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__or2b_1 _15840_ (.A(_08479_),
    .B_N(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__xnor2_1 _15841_ (.A(_08137_),
    .B(_08143_),
    .Y(_08486_));
 sky130_fd_sc_hd__a21o_1 _15842_ (.A1(_08478_),
    .A2(_08485_),
    .B1(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__nand3_1 _15843_ (.A(_08478_),
    .B(_08485_),
    .C(_08486_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand2_1 _15844_ (.A(_08487_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__nand2_1 _15845_ (.A(_07945_),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .Y(_08490_));
 sky130_fd_sc_hd__and2_4 _15846_ (.A(_08124_),
    .B(_08490_),
    .X(_08491_));
 sky130_fd_sc_hd__or4_4 _15847_ (.A(_08129_),
    .B(_08047_),
    .C(_08135_),
    .D(_08491_),
    .X(_08492_));
 sky130_fd_sc_hd__buf_4 _15848_ (.A(_08129_),
    .X(_08493_));
 sky130_fd_sc_hd__o22ai_4 _15849_ (.A1(_08047_),
    .A2(_08135_),
    .B1(_08491_),
    .B2(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__o21bai_1 _15850_ (.A1(_08113_),
    .A2(_08139_),
    .B1_N(_08140_),
    .Y(_08495_));
 sky130_fd_sc_hd__xnor2_1 _15851_ (.A(_08495_),
    .B(_08141_),
    .Y(_08496_));
 sky130_fd_sc_hd__nor2_1 _15852_ (.A(_08097_),
    .B(_08491_),
    .Y(_08497_));
 sky130_fd_sc_hd__or2_1 _15853_ (.A(_08074_),
    .B(_08125_),
    .X(_08498_));
 sky130_fd_sc_hd__or3_1 _15854_ (.A(_08084_),
    .B(_08041_),
    .C(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__o22ai_1 _15855_ (.A1(_08109_),
    .A2(_08042_),
    .B1(_08125_),
    .B2(_08084_),
    .Y(_08500_));
 sky130_fd_sc_hd__and2_1 _15856_ (.A(_08499_),
    .B(_08500_),
    .X(_08501_));
 sky130_fd_sc_hd__a21boi_1 _15857_ (.A1(_08497_),
    .A2(_08501_),
    .B1_N(_08499_),
    .Y(_08502_));
 sky130_fd_sc_hd__xor2_1 _15858_ (.A(_08496_),
    .B(_08502_),
    .X(_08503_));
 sky130_fd_sc_hd__nor2_1 _15859_ (.A(_08496_),
    .B(_08502_),
    .Y(_08504_));
 sky130_fd_sc_hd__a31o_1 _15860_ (.A1(_08492_),
    .A2(_08494_),
    .A3(_08503_),
    .B1(_08504_),
    .X(_08505_));
 sky130_fd_sc_hd__or2b_1 _15861_ (.A(_08489_),
    .B_N(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__nand2_1 _15862_ (.A(_08152_),
    .B(_08153_),
    .Y(_08507_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_08154_),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__a21oi_4 _15864_ (.A1(_08487_),
    .A2(_08506_),
    .B1(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__and2b_1 _15865_ (.A_N(_08467_),
    .B(_08464_),
    .X(_08510_));
 sky130_fd_sc_hd__xnor2_4 _15866_ (.A(_08510_),
    .B(_08466_),
    .Y(_08511_));
 sky130_fd_sc_hd__xnor2_1 _15867_ (.A(_08460_),
    .B(_08461_),
    .Y(_08512_));
 sky130_fd_sc_hd__xnor2_1 _15868_ (.A(_08456_),
    .B(_08457_),
    .Y(_08513_));
 sky130_fd_sc_hd__xnor2_2 _15869_ (.A(_08451_),
    .B(_08453_),
    .Y(_08514_));
 sky130_fd_sc_hd__and2_1 _15870_ (.A(\rbzero.wall_tracer.visualWallDist[-12] ),
    .B(_07925_),
    .X(_08515_));
 sky130_fd_sc_hd__and3_1 _15871_ (.A(_08199_),
    .B(_08201_),
    .C(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__xor2_2 _15872_ (.A(_08448_),
    .B(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__or2_1 _15873_ (.A(_05195_),
    .B(_08226_),
    .X(_08518_));
 sky130_fd_sc_hd__buf_4 _15874_ (.A(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__nor2_1 _15875_ (.A(_07974_),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__and4_1 _15876_ (.A(_07601_),
    .B(_04014_),
    .C(_05197_),
    .D(_07992_),
    .X(_08521_));
 sky130_fd_sc_hd__xnor2_1 _15877_ (.A(_08520_),
    .B(_08521_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand2_1 _15878_ (.A(_08445_),
    .B(_08250_),
    .Y(_08523_));
 sky130_fd_sc_hd__and2_1 _15879_ (.A(_08520_),
    .B(_08521_),
    .X(_08524_));
 sky130_fd_sc_hd__o21ba_1 _15880_ (.A1(_08522_),
    .A2(_08523_),
    .B1_N(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__xor2_2 _15881_ (.A(_08517_),
    .B(_08525_),
    .X(_08526_));
 sky130_fd_sc_hd__nand2_1 _15882_ (.A(_08476_),
    .B(_08473_),
    .Y(_08527_));
 sky130_fd_sc_hd__xnor2_2 _15883_ (.A(_08527_),
    .B(_08474_),
    .Y(_08528_));
 sky130_fd_sc_hd__nor2_1 _15884_ (.A(_08517_),
    .B(_08525_),
    .Y(_08529_));
 sky130_fd_sc_hd__a21oi_2 _15885_ (.A1(_08526_),
    .A2(_08528_),
    .B1(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__xor2_2 _15886_ (.A(_08514_),
    .B(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__xnor2_2 _15887_ (.A(_08484_),
    .B(_08479_),
    .Y(_08532_));
 sky130_fd_sc_hd__nor2_1 _15888_ (.A(_08514_),
    .B(_08530_),
    .Y(_08533_));
 sky130_fd_sc_hd__a21oi_1 _15889_ (.A1(_08531_),
    .A2(_08532_),
    .B1(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__xor2_1 _15890_ (.A(_08513_),
    .B(_08534_),
    .X(_08535_));
 sky130_fd_sc_hd__xnor2_1 _15891_ (.A(_08505_),
    .B(_08489_),
    .Y(_08536_));
 sky130_fd_sc_hd__nor2_1 _15892_ (.A(_08513_),
    .B(_08534_),
    .Y(_08537_));
 sky130_fd_sc_hd__a21oi_1 _15893_ (.A1(_08535_),
    .A2(_08536_),
    .B1(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__xor2_1 _15894_ (.A(_08512_),
    .B(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__and3_1 _15895_ (.A(_08487_),
    .B(_08506_),
    .C(_08508_),
    .X(_08540_));
 sky130_fd_sc_hd__nor2_1 _15896_ (.A(_08509_),
    .B(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__nor2_1 _15897_ (.A(_08512_),
    .B(_08538_),
    .Y(_08542_));
 sky130_fd_sc_hd__a21oi_2 _15898_ (.A1(_08539_),
    .A2(_08541_),
    .B1(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__xor2_4 _15899_ (.A(_08511_),
    .B(_08543_),
    .X(_08544_));
 sky130_fd_sc_hd__nor2_1 _15900_ (.A(_08511_),
    .B(_08543_),
    .Y(_08545_));
 sky130_fd_sc_hd__a21oi_2 _15901_ (.A1(_08509_),
    .A2(_08544_),
    .B1(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__nor2_2 _15902_ (.A(_08470_),
    .B(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__and2_1 _15903_ (.A(_08470_),
    .B(_08546_),
    .X(_08548_));
 sky130_fd_sc_hd__nor2_4 _15904_ (.A(_08547_),
    .B(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__xnor2_4 _15905_ (.A(_08509_),
    .B(_08544_),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2_1 _15906_ (.A(_08483_),
    .B(_08480_),
    .Y(_08551_));
 sky130_fd_sc_hd__xor2_1 _15907_ (.A(_08551_),
    .B(_08481_),
    .X(_08552_));
 sky130_fd_sc_hd__or3_1 _15908_ (.A(_07988_),
    .B(_07938_),
    .C(_07939_),
    .X(_08553_));
 sky130_fd_sc_hd__xor2_1 _15909_ (.A(_08475_),
    .B(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__nor2_1 _15910_ (.A(_08008_),
    .B(_07967_),
    .Y(_08555_));
 sky130_fd_sc_hd__a2bb2o_1 _15911_ (.A1_N(_08475_),
    .A2_N(_08553_),
    .B1(_08554_),
    .B2(_08555_),
    .X(_08556_));
 sky130_fd_sc_hd__or2b_1 _15912_ (.A(_08552_),
    .B_N(_08556_),
    .X(_08557_));
 sky130_fd_sc_hd__xor2_1 _15913_ (.A(_08556_),
    .B(_08552_),
    .X(_08558_));
 sky130_fd_sc_hd__or3_1 _15914_ (.A(_07923_),
    .B(_08102_),
    .C(_08103_),
    .X(_08559_));
 sky130_fd_sc_hd__nor2_1 _15915_ (.A(_07959_),
    .B(_08042_),
    .Y(_08560_));
 sky130_fd_sc_hd__xor2_1 _15916_ (.A(_08482_),
    .B(_08559_),
    .X(_08561_));
 sky130_fd_sc_hd__a2bb2o_1 _15917_ (.A1_N(_08482_),
    .A2_N(_08559_),
    .B1(_08560_),
    .B2(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__or2b_1 _15918_ (.A(_08558_),
    .B_N(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__nand2_1 _15919_ (.A(_08492_),
    .B(_08494_),
    .Y(_08564_));
 sky130_fd_sc_hd__xor2_1 _15920_ (.A(_08564_),
    .B(_08503_),
    .X(_08565_));
 sky130_fd_sc_hd__a21o_1 _15921_ (.A1(_08557_),
    .A2(_08563_),
    .B1(_08565_),
    .X(_08566_));
 sky130_fd_sc_hd__nand3_1 _15922_ (.A(_08557_),
    .B(_08563_),
    .C(_08565_),
    .Y(_08567_));
 sky130_fd_sc_hd__nand2_1 _15923_ (.A(_08566_),
    .B(_08567_),
    .Y(_08568_));
 sky130_fd_sc_hd__xnor2_2 _15924_ (.A(_08497_),
    .B(_08501_),
    .Y(_08569_));
 sky130_fd_sc_hd__buf_4 _15925_ (.A(_08084_),
    .X(_08570_));
 sky130_fd_sc_hd__or2_1 _15926_ (.A(_08109_),
    .B(_08491_),
    .X(_08571_));
 sky130_fd_sc_hd__a21boi_4 _15927_ (.A1(_07945_),
    .A2(\rbzero.wall_tracer.stepDistX[-12] ),
    .B1_N(_08135_),
    .Y(_08572_));
 sky130_fd_sc_hd__or2_1 _15928_ (.A(_08096_),
    .B(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__a21oi_1 _15929_ (.A1(_08124_),
    .A2(_08490_),
    .B1(_08084_),
    .Y(_08574_));
 sky130_fd_sc_hd__xnor2_1 _15930_ (.A(_08498_),
    .B(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__or2b_1 _15931_ (.A(_08573_),
    .B_N(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__o31a_1 _15932_ (.A1(_08570_),
    .A2(_08128_),
    .A3(_08571_),
    .B1(_08576_),
    .X(_08577_));
 sky130_fd_sc_hd__xnor2_2 _15933_ (.A(_08569_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__buf_2 _15934_ (.A(_08572_),
    .X(_08579_));
 sky130_fd_sc_hd__or2_2 _15935_ (.A(_08129_),
    .B(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__or2_1 _15936_ (.A(_08569_),
    .B(_08577_),
    .X(_08581_));
 sky130_fd_sc_hd__o21ai_2 _15937_ (.A1(_08578_),
    .A2(_08580_),
    .B1(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__or2b_1 _15938_ (.A(_08568_),
    .B_N(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__a21oi_4 _15939_ (.A1(_08566_),
    .A2(_08583_),
    .B1(_08492_),
    .Y(_08584_));
 sky130_fd_sc_hd__xnor2_1 _15940_ (.A(_08539_),
    .B(_08541_),
    .Y(_08585_));
 sky130_fd_sc_hd__xnor2_1 _15941_ (.A(_08535_),
    .B(_08536_),
    .Y(_08586_));
 sky130_fd_sc_hd__xnor2_2 _15942_ (.A(_08531_),
    .B(_08532_),
    .Y(_08587_));
 sky130_fd_sc_hd__xnor2_2 _15943_ (.A(_08526_),
    .B(_08528_),
    .Y(_08588_));
 sky130_fd_sc_hd__xor2_2 _15944_ (.A(_08555_),
    .B(_08554_),
    .X(_08589_));
 sky130_fd_sc_hd__xnor2_1 _15945_ (.A(_08522_),
    .B(_08523_),
    .Y(_08590_));
 sky130_fd_sc_hd__and4_1 _15946_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_04014_),
    .C(_05197_),
    .D(_07992_),
    .X(_08591_));
 sky130_fd_sc_hd__and4_1 _15947_ (.A(_07601_),
    .B(_04014_),
    .C(_07990_),
    .D(_07927_),
    .X(_08592_));
 sky130_fd_sc_hd__xnor2_1 _15948_ (.A(_08591_),
    .B(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_2 _15949_ (.A(_07990_),
    .B(_08515_),
    .Y(_08594_));
 sky130_fd_sc_hd__or2_1 _15950_ (.A(_07974_),
    .B(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__nand2_1 _15951_ (.A(_08591_),
    .B(_08592_),
    .Y(_08596_));
 sky130_fd_sc_hd__o21a_1 _15952_ (.A1(_08593_),
    .A2(_08595_),
    .B1(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__xor2_1 _15953_ (.A(_08590_),
    .B(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__nor2_1 _15954_ (.A(_08590_),
    .B(_08597_),
    .Y(_08599_));
 sky130_fd_sc_hd__a21oi_2 _15955_ (.A1(_08589_),
    .A2(_08598_),
    .B1(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__xor2_2 _15956_ (.A(_08588_),
    .B(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__xnor2_2 _15957_ (.A(_08562_),
    .B(_08558_),
    .Y(_08602_));
 sky130_fd_sc_hd__nor2_1 _15958_ (.A(_08588_),
    .B(_08600_),
    .Y(_08603_));
 sky130_fd_sc_hd__a21oi_2 _15959_ (.A1(_08601_),
    .A2(_08602_),
    .B1(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__xor2_2 _15960_ (.A(_08587_),
    .B(_08604_),
    .X(_08605_));
 sky130_fd_sc_hd__xnor2_2 _15961_ (.A(_08582_),
    .B(_08568_),
    .Y(_08606_));
 sky130_fd_sc_hd__nor2_1 _15962_ (.A(_08587_),
    .B(_08604_),
    .Y(_08607_));
 sky130_fd_sc_hd__a21oi_1 _15963_ (.A1(_08605_),
    .A2(_08606_),
    .B1(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__xor2_1 _15964_ (.A(_08586_),
    .B(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__and3_1 _15965_ (.A(_08492_),
    .B(_08566_),
    .C(_08583_),
    .X(_08610_));
 sky130_fd_sc_hd__nor2_1 _15966_ (.A(_08584_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__nor2_1 _15967_ (.A(_08586_),
    .B(_08608_),
    .Y(_08612_));
 sky130_fd_sc_hd__a21oi_1 _15968_ (.A1(_08609_),
    .A2(_08611_),
    .B1(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand2_1 _15969_ (.A(_08585_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__nor2_1 _15970_ (.A(_08585_),
    .B(_08613_),
    .Y(_08615_));
 sky130_fd_sc_hd__a21oi_4 _15971_ (.A1(_08584_),
    .A2(_08614_),
    .B1(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__xor2_2 _15972_ (.A(_08550_),
    .B(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__and2b_1 _15973_ (.A_N(_08615_),
    .B(_08614_),
    .X(_08618_));
 sky130_fd_sc_hd__xnor2_4 _15974_ (.A(_08584_),
    .B(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__xnor2_1 _15975_ (.A(_08609_),
    .B(_08611_),
    .Y(_08620_));
 sky130_fd_sc_hd__xnor2_2 _15976_ (.A(_08605_),
    .B(_08606_),
    .Y(_08621_));
 sky130_fd_sc_hd__xnor2_2 _15977_ (.A(_08601_),
    .B(_08602_),
    .Y(_08622_));
 sky130_fd_sc_hd__or3b_2 _15978_ (.A(_07912_),
    .B(_08328_),
    .C_N(_08040_),
    .X(_08623_));
 sky130_fd_sc_hd__nor2_1 _15979_ (.A(_07958_),
    .B(_08128_),
    .Y(_08624_));
 sky130_fd_sc_hd__or3_1 _15980_ (.A(_07912_),
    .B(_08102_),
    .C(_08103_),
    .X(_08625_));
 sky130_fd_sc_hd__inv_2 _15981_ (.A(_07923_),
    .Y(_08626_));
 sky130_fd_sc_hd__and3_1 _15982_ (.A(_08626_),
    .B(_08039_),
    .C(_08040_),
    .X(_08627_));
 sky130_fd_sc_hd__xnor2_1 _15983_ (.A(_08625_),
    .B(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__a2bb2o_1 _15984_ (.A1_N(_08559_),
    .A2_N(_08623_),
    .B1(_08624_),
    .B2(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__or3_1 _15985_ (.A(_07980_),
    .B(_07938_),
    .C(_07939_),
    .X(_08630_));
 sky130_fd_sc_hd__or3_1 _15986_ (.A(_07988_),
    .B(_07964_),
    .C(_07965_),
    .X(_08631_));
 sky130_fd_sc_hd__xor2_1 _15987_ (.A(_08630_),
    .B(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__nor2_1 _15988_ (.A(_08008_),
    .B(_08022_),
    .Y(_08633_));
 sky130_fd_sc_hd__a2bb2o_1 _15989_ (.A1_N(_08630_),
    .A2_N(_08631_),
    .B1(_08632_),
    .B2(_08633_),
    .X(_08634_));
 sky130_fd_sc_hd__or2_1 _15990_ (.A(_07958_),
    .B(_08041_),
    .X(_08635_));
 sky130_fd_sc_hd__xnor2_1 _15991_ (.A(_08635_),
    .B(_08561_),
    .Y(_08636_));
 sky130_fd_sc_hd__xnor2_1 _15992_ (.A(_08634_),
    .B(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__xnor2_1 _15993_ (.A(_08629_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__xnor2_1 _15994_ (.A(_08589_),
    .B(_08598_),
    .Y(_08639_));
 sky130_fd_sc_hd__xor2_1 _15995_ (.A(_08633_),
    .B(_08632_),
    .X(_08640_));
 sky130_fd_sc_hd__xnor2_1 _15996_ (.A(_08593_),
    .B(_08595_),
    .Y(_08641_));
 sky130_fd_sc_hd__or4b_2 _15997_ (.A(_07598_),
    .B(_07951_),
    .C(_05207_),
    .D_N(_07927_),
    .X(_08642_));
 sky130_fd_sc_hd__and4_1 _15998_ (.A(_07601_),
    .B(_04014_),
    .C(_07990_),
    .D(_07936_),
    .X(_08643_));
 sky130_fd_sc_hd__xnor2_2 _15999_ (.A(_08642_),
    .B(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__nor2_1 _16000_ (.A(_07994_),
    .B(_08594_),
    .Y(_08645_));
 sky130_fd_sc_hd__and2b_1 _16001_ (.A_N(_08642_),
    .B(_08643_),
    .X(_08646_));
 sky130_fd_sc_hd__a21oi_1 _16002_ (.A1(_08644_),
    .A2(_08645_),
    .B1(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__xor2_1 _16003_ (.A(_08641_),
    .B(_08647_),
    .X(_08648_));
 sky130_fd_sc_hd__nor2_1 _16004_ (.A(_08641_),
    .B(_08647_),
    .Y(_08649_));
 sky130_fd_sc_hd__a21oi_1 _16005_ (.A1(_08640_),
    .A2(_08648_),
    .B1(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__xor2_1 _16006_ (.A(_08639_),
    .B(_08650_),
    .X(_08651_));
 sky130_fd_sc_hd__nor2_1 _16007_ (.A(_08639_),
    .B(_08650_),
    .Y(_08652_));
 sky130_fd_sc_hd__a21oi_2 _16008_ (.A1(_08638_),
    .A2(_08651_),
    .B1(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__xor2_2 _16009_ (.A(_08622_),
    .B(_08653_),
    .X(_08654_));
 sky130_fd_sc_hd__or2b_1 _16010_ (.A(_08637_),
    .B_N(_08629_),
    .X(_08655_));
 sky130_fd_sc_hd__a21bo_1 _16011_ (.A1(_08634_),
    .A2(_08636_),
    .B1_N(_08655_),
    .X(_08656_));
 sky130_fd_sc_hd__xnor2_2 _16012_ (.A(_08578_),
    .B(_08580_),
    .Y(_08657_));
 sky130_fd_sc_hd__xor2_2 _16013_ (.A(_08656_),
    .B(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__xnor2_1 _16014_ (.A(_08573_),
    .B(_08575_),
    .Y(_08659_));
 sky130_fd_sc_hd__nor2_1 _16015_ (.A(_08111_),
    .B(_08579_),
    .Y(_08660_));
 sky130_fd_sc_hd__and2_1 _16016_ (.A(_08574_),
    .B(_08660_),
    .X(_08661_));
 sky130_fd_sc_hd__nand2_1 _16017_ (.A(_08659_),
    .B(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__xor2_2 _16018_ (.A(_08658_),
    .B(_08662_),
    .X(_08663_));
 sky130_fd_sc_hd__nor2_1 _16019_ (.A(_08622_),
    .B(_08653_),
    .Y(_08664_));
 sky130_fd_sc_hd__a21oi_1 _16020_ (.A1(_08654_),
    .A2(_08663_),
    .B1(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__xnor2_2 _16021_ (.A(_08621_),
    .B(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__or2b_1 _16022_ (.A(_08657_),
    .B_N(_08656_),
    .X(_08667_));
 sky130_fd_sc_hd__o21a_2 _16023_ (.A1(_08658_),
    .A2(_08662_),
    .B1(_08667_),
    .X(_08668_));
 sky130_fd_sc_hd__or2_1 _16024_ (.A(_08621_),
    .B(_08665_),
    .X(_08669_));
 sky130_fd_sc_hd__o21a_1 _16025_ (.A1(_08666_),
    .A2(_08668_),
    .B1(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__nor2_1 _16026_ (.A(_08620_),
    .B(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__and2b_1 _16027_ (.A_N(_08619_),
    .B(_08671_),
    .X(_08672_));
 sky130_fd_sc_hd__nor2_1 _16028_ (.A(_08617_),
    .B(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__clkbuf_4 _16029_ (.A(_08019_),
    .X(_08674_));
 sky130_fd_sc_hd__or3_2 _16030_ (.A(_07980_),
    .B(_08674_),
    .C(_08020_),
    .X(_08675_));
 sky130_fd_sc_hd__or3_1 _16031_ (.A(_07980_),
    .B(_07964_),
    .C(_07965_),
    .X(_08676_));
 sky130_fd_sc_hd__or3_1 _16032_ (.A(_07988_),
    .B(_08674_),
    .C(_08020_),
    .X(_08677_));
 sky130_fd_sc_hd__and2_1 _16033_ (.A(_08676_),
    .B(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__or2_1 _16034_ (.A(_08008_),
    .B(_08104_),
    .X(_08679_));
 sky130_fd_sc_hd__o22a_1 _16035_ (.A1(_08631_),
    .A2(_08675_),
    .B1(_08678_),
    .B2(_08679_),
    .X(_08680_));
 sky130_fd_sc_hd__xnor2_1 _16036_ (.A(_08624_),
    .B(_08628_),
    .Y(_08681_));
 sky130_fd_sc_hd__or2_1 _16037_ (.A(_08680_),
    .B(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__xnor2_1 _16038_ (.A(_08680_),
    .B(_08681_),
    .Y(_08683_));
 sky130_fd_sc_hd__or2_1 _16039_ (.A(_07958_),
    .B(_08491_),
    .X(_08684_));
 sky130_fd_sc_hd__nor2_1 _16040_ (.A(_07923_),
    .B(_08125_),
    .Y(_08685_));
 sky130_fd_sc_hd__xnor2_1 _16041_ (.A(_08623_),
    .B(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__or2b_1 _16042_ (.A(_08684_),
    .B_N(_08686_),
    .X(_08687_));
 sky130_fd_sc_hd__o31ai_2 _16043_ (.A1(_08284_),
    .A2(_08128_),
    .A3(_08623_),
    .B1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__or2b_1 _16044_ (.A(_08683_),
    .B_N(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__or2_1 _16045_ (.A(_08659_),
    .B(_08661_),
    .X(_08690_));
 sky130_fd_sc_hd__nand2_1 _16046_ (.A(_08662_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__a21oi_4 _16047_ (.A1(_08682_),
    .A2(_08689_),
    .B1(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__xnor2_2 _16048_ (.A(_08654_),
    .B(_08663_),
    .Y(_08693_));
 sky130_fd_sc_hd__and3_1 _16049_ (.A(_08682_),
    .B(_08689_),
    .C(_08691_),
    .X(_08694_));
 sky130_fd_sc_hd__nor2_2 _16050_ (.A(_08692_),
    .B(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__xnor2_1 _16051_ (.A(_08638_),
    .B(_08651_),
    .Y(_08696_));
 sky130_fd_sc_hd__xnor2_1 _16052_ (.A(_08688_),
    .B(_08683_),
    .Y(_08697_));
 sky130_fd_sc_hd__xnor2_1 _16053_ (.A(_08640_),
    .B(_08648_),
    .Y(_08698_));
 sky130_fd_sc_hd__xor2_1 _16054_ (.A(_08676_),
    .B(_08677_),
    .X(_08699_));
 sky130_fd_sc_hd__xnor2_2 _16055_ (.A(_08679_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__xnor2_2 _16056_ (.A(_08644_),
    .B(_08645_),
    .Y(_08701_));
 sky130_fd_sc_hd__and4_1 _16057_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_04014_),
    .C(_07990_),
    .D(_07936_),
    .X(_08702_));
 sky130_fd_sc_hd__and4_1 _16058_ (.A(_07601_),
    .B(_08148_),
    .C(_07990_),
    .D(_07962_),
    .X(_08703_));
 sky130_fd_sc_hd__xor2_2 _16059_ (.A(_08702_),
    .B(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__buf_4 _16060_ (.A(_07929_),
    .X(_08705_));
 sky130_fd_sc_hd__nor2_1 _16061_ (.A(_08594_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__and2_1 _16062_ (.A(_08702_),
    .B(_08703_),
    .X(_08707_));
 sky130_fd_sc_hd__a21oi_2 _16063_ (.A1(_08704_),
    .A2(_08706_),
    .B1(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__xor2_2 _16064_ (.A(_08701_),
    .B(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__nor2_1 _16065_ (.A(_08701_),
    .B(_08708_),
    .Y(_08710_));
 sky130_fd_sc_hd__a21o_1 _16066_ (.A1(_08700_),
    .A2(_08709_),
    .B1(_08710_),
    .X(_08711_));
 sky130_fd_sc_hd__xnor2_1 _16067_ (.A(_08698_),
    .B(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__and2b_1 _16068_ (.A_N(_08698_),
    .B(_08711_),
    .X(_08713_));
 sky130_fd_sc_hd__a21oi_1 _16069_ (.A1(_08697_),
    .A2(_08712_),
    .B1(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_1 _16070_ (.A(_08696_),
    .B(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__nor2_1 _16071_ (.A(_08696_),
    .B(_08714_),
    .Y(_08716_));
 sky130_fd_sc_hd__a21oi_2 _16072_ (.A1(_08695_),
    .A2(_08715_),
    .B1(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__xor2_2 _16073_ (.A(_08693_),
    .B(_08717_),
    .X(_08718_));
 sky130_fd_sc_hd__xnor2_2 _16074_ (.A(_08692_),
    .B(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__or3_2 _16075_ (.A(_07989_),
    .B(_08102_),
    .C(_08103_),
    .X(_08720_));
 sky130_fd_sc_hd__xor2_1 _16076_ (.A(_08675_),
    .B(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__nor2_1 _16077_ (.A(_08008_),
    .B(_08042_),
    .Y(_08722_));
 sky130_fd_sc_hd__a2bb2o_1 _16078_ (.A1_N(_08675_),
    .A2_N(_08720_),
    .B1(_08721_),
    .B2(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__xnor2_1 _16079_ (.A(_08684_),
    .B(_08686_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand2_1 _16080_ (.A(_08723_),
    .B(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__xnor2_1 _16081_ (.A(_08723_),
    .B(_08724_),
    .Y(_08726_));
 sky130_fd_sc_hd__or2_1 _16082_ (.A(_08283_),
    .B(_08491_),
    .X(_08727_));
 sky130_fd_sc_hd__or2_1 _16083_ (.A(_07958_),
    .B(_08572_),
    .X(_08728_));
 sky130_fd_sc_hd__or2_1 _16084_ (.A(_07912_),
    .B(_08125_),
    .X(_08729_));
 sky130_fd_sc_hd__a21oi_1 _16085_ (.A1(_08124_),
    .A2(_08490_),
    .B1(_07924_),
    .Y(_08730_));
 sky130_fd_sc_hd__xnor2_1 _16086_ (.A(_08729_),
    .B(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__or2b_1 _16087_ (.A(_08728_),
    .B_N(_08731_),
    .X(_08732_));
 sky130_fd_sc_hd__o31ai_2 _16088_ (.A1(_08284_),
    .A2(_08128_),
    .A3(_08727_),
    .B1(_08732_),
    .Y(_08733_));
 sky130_fd_sc_hd__or2b_1 _16089_ (.A(_08726_),
    .B_N(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__o21a_1 _16090_ (.A1(_08570_),
    .A2(_08579_),
    .B1(_08571_),
    .X(_08735_));
 sky130_fd_sc_hd__or2_1 _16091_ (.A(_08661_),
    .B(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__a21oi_2 _16092_ (.A1(_08725_),
    .A2(_08734_),
    .B1(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__and2b_1 _16093_ (.A_N(_08716_),
    .B(_08715_),
    .X(_08738_));
 sky130_fd_sc_hd__xnor2_2 _16094_ (.A(_08695_),
    .B(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__xnor2_1 _16095_ (.A(_08697_),
    .B(_08712_),
    .Y(_08740_));
 sky130_fd_sc_hd__xnor2_1 _16096_ (.A(_08733_),
    .B(_08726_),
    .Y(_08741_));
 sky130_fd_sc_hd__xnor2_2 _16097_ (.A(_08700_),
    .B(_08709_),
    .Y(_08742_));
 sky130_fd_sc_hd__xor2_1 _16098_ (.A(_08722_),
    .B(_08721_),
    .X(_08743_));
 sky130_fd_sc_hd__xnor2_2 _16099_ (.A(_08704_),
    .B(_08706_),
    .Y(_08744_));
 sky130_fd_sc_hd__o22ai_2 _16100_ (.A1(_08519_),
    .A2(_08075_),
    .B1(_08674_),
    .B2(_08377_),
    .Y(_08745_));
 sky130_fd_sc_hd__nor2_1 _16101_ (.A(_08594_),
    .B(_07938_),
    .Y(_08746_));
 sky130_fd_sc_hd__nand2_2 _16102_ (.A(_07601_),
    .B(_08227_),
    .Y(_08747_));
 sky130_fd_sc_hd__or3_1 _16103_ (.A(_07964_),
    .B(_08674_),
    .C(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__a21boi_2 _16104_ (.A1(_08745_),
    .A2(_08746_),
    .B1_N(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__xor2_1 _16105_ (.A(_08744_),
    .B(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__nor2_1 _16106_ (.A(_08744_),
    .B(_08749_),
    .Y(_08751_));
 sky130_fd_sc_hd__a21oi_1 _16107_ (.A1(_08743_),
    .A2(_08750_),
    .B1(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__xor2_1 _16108_ (.A(_08742_),
    .B(_08752_),
    .X(_08753_));
 sky130_fd_sc_hd__nor2_1 _16109_ (.A(_08742_),
    .B(_08752_),
    .Y(_08754_));
 sky130_fd_sc_hd__a21oi_1 _16110_ (.A1(_08741_),
    .A2(_08753_),
    .B1(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(_08740_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__and3_1 _16112_ (.A(_08725_),
    .B(_08734_),
    .C(_08736_),
    .X(_08757_));
 sky130_fd_sc_hd__nor2_1 _16113_ (.A(_08737_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__nor2_1 _16114_ (.A(_08740_),
    .B(_08755_),
    .Y(_08759_));
 sky130_fd_sc_hd__a21oi_2 _16115_ (.A1(_08756_),
    .A2(_08758_),
    .B1(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__xor2_2 _16116_ (.A(_08739_),
    .B(_08760_),
    .X(_08761_));
 sky130_fd_sc_hd__nor2_1 _16117_ (.A(_08739_),
    .B(_08760_),
    .Y(_08762_));
 sky130_fd_sc_hd__a21oi_2 _16118_ (.A1(_08737_),
    .A2(_08761_),
    .B1(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__xor2_2 _16119_ (.A(_08719_),
    .B(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__and2b_1 _16120_ (.A_N(_08759_),
    .B(_08756_),
    .X(_08765_));
 sky130_fd_sc_hd__xnor2_1 _16121_ (.A(_08765_),
    .B(_08758_),
    .Y(_08766_));
 sky130_fd_sc_hd__buf_4 _16122_ (.A(_08284_),
    .X(_08767_));
 sky130_fd_sc_hd__or2_1 _16123_ (.A(_08008_),
    .B(_08128_),
    .X(_08768_));
 sky130_fd_sc_hd__or3_1 _16124_ (.A(_07980_),
    .B(_08102_),
    .C(_08103_),
    .X(_08769_));
 sky130_fd_sc_hd__o21a_1 _16125_ (.A1(_08180_),
    .A2(_08042_),
    .B1(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__or3_1 _16126_ (.A(_07981_),
    .B(_08042_),
    .C(_08720_),
    .X(_08771_));
 sky130_fd_sc_hd__o21a_1 _16127_ (.A1(_08768_),
    .A2(_08770_),
    .B1(_08771_),
    .X(_08772_));
 sky130_fd_sc_hd__xnor2_1 _16128_ (.A(_08728_),
    .B(_08731_),
    .Y(_08773_));
 sky130_fd_sc_hd__or2b_1 _16129_ (.A(_08772_),
    .B_N(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__or2b_1 _16130_ (.A(_08773_),
    .B_N(_08772_),
    .X(_08775_));
 sky130_fd_sc_hd__nand2_1 _16131_ (.A(_08774_),
    .B(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__o41a_1 _16132_ (.A1(_08767_),
    .A2(_08579_),
    .A3(_08727_),
    .A4(_08776_),
    .B1(_08774_),
    .X(_08777_));
 sky130_fd_sc_hd__xnor2_1 _16133_ (.A(_08660_),
    .B(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__xnor2_1 _16134_ (.A(_08741_),
    .B(_08753_),
    .Y(_08779_));
 sky130_fd_sc_hd__nand2_1 _16135_ (.A(_08743_),
    .B(_08750_),
    .Y(_08780_));
 sky130_fd_sc_hd__or2_1 _16136_ (.A(_08743_),
    .B(_08750_),
    .X(_08781_));
 sky130_fd_sc_hd__and3_1 _16137_ (.A(_08748_),
    .B(_08745_),
    .C(_08746_),
    .X(_08782_));
 sky130_fd_sc_hd__a21oi_1 _16138_ (.A1(_08748_),
    .A2(_08745_),
    .B1(_08746_),
    .Y(_08783_));
 sky130_fd_sc_hd__o22a_1 _16139_ (.A1(_08519_),
    .A2(_08674_),
    .B1(_08112_),
    .B2(_08377_),
    .X(_08784_));
 sky130_fd_sc_hd__or3_1 _16140_ (.A(_08674_),
    .B(_08112_),
    .C(_08747_),
    .X(_08785_));
 sky130_fd_sc_hd__o31a_1 _16141_ (.A1(_08594_),
    .A2(_08075_),
    .A3(_08784_),
    .B1(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__o21ai_2 _16142_ (.A1(_08782_),
    .A2(_08783_),
    .B1(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__and3_1 _16143_ (.A(_08266_),
    .B(_08039_),
    .C(_08040_),
    .X(_08788_));
 sky130_fd_sc_hd__xnor2_1 _16144_ (.A(_08769_),
    .B(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__xnor2_1 _16145_ (.A(_08768_),
    .B(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__or3_1 _16146_ (.A(_08782_),
    .B(_08783_),
    .C(_08786_),
    .X(_08791_));
 sky130_fd_sc_hd__a21bo_1 _16147_ (.A1(_08787_),
    .A2(_08790_),
    .B1_N(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__nor3_1 _16148_ (.A(_08284_),
    .B(_08579_),
    .C(_08727_),
    .Y(_08793_));
 sky130_fd_sc_hd__xnor2_1 _16149_ (.A(_08776_),
    .B(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_1 _16150_ (.A(_08780_),
    .B(_08781_),
    .Y(_08795_));
 sky130_fd_sc_hd__xnor2_1 _16151_ (.A(_08795_),
    .B(_08792_),
    .Y(_08796_));
 sky130_fd_sc_hd__a32oi_2 _16152_ (.A1(_08780_),
    .A2(_08781_),
    .A3(_08792_),
    .B1(_08794_),
    .B2(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__nand2_1 _16153_ (.A(_08779_),
    .B(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__nor2_1 _16154_ (.A(_08779_),
    .B(_08797_),
    .Y(_08799_));
 sky130_fd_sc_hd__a21oi_1 _16155_ (.A1(_08778_),
    .A2(_08798_),
    .B1(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__or2_1 _16156_ (.A(_08766_),
    .B(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__buf_4 _16157_ (.A(_08111_),
    .X(_08802_));
 sky130_fd_sc_hd__or3_1 _16158_ (.A(_08802_),
    .B(_08579_),
    .C(_08777_),
    .X(_08803_));
 sky130_fd_sc_hd__xnor2_1 _16159_ (.A(_08766_),
    .B(_08800_),
    .Y(_08804_));
 sky130_fd_sc_hd__or2_1 _16160_ (.A(_08803_),
    .B(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__xnor2_2 _16161_ (.A(_08737_),
    .B(_08761_),
    .Y(_08806_));
 sky130_fd_sc_hd__a21oi_4 _16162_ (.A1(_08801_),
    .A2(_08805_),
    .B1(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__xnor2_4 _16163_ (.A(_08666_),
    .B(_08668_),
    .Y(_08808_));
 sky130_fd_sc_hd__nor2_1 _16164_ (.A(_08693_),
    .B(_08717_),
    .Y(_08809_));
 sky130_fd_sc_hd__a21oi_2 _16165_ (.A1(_08692_),
    .A2(_08718_),
    .B1(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__xor2_4 _16166_ (.A(_08808_),
    .B(_08810_),
    .X(_08811_));
 sky130_fd_sc_hd__xnor2_1 _16167_ (.A(_08794_),
    .B(_08796_),
    .Y(_08812_));
 sky130_fd_sc_hd__and3_1 _16168_ (.A(_08791_),
    .B(_08787_),
    .C(_08790_),
    .X(_08813_));
 sky130_fd_sc_hd__a21oi_1 _16169_ (.A1(_08791_),
    .A2(_08787_),
    .B1(_08790_),
    .Y(_08814_));
 sky130_fd_sc_hd__or2_1 _16170_ (.A(_08813_),
    .B(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__clkbuf_4 _16171_ (.A(_08594_),
    .X(_08816_));
 sky130_fd_sc_hd__nor3_1 _16172_ (.A(_08674_),
    .B(_08112_),
    .C(_08747_),
    .Y(_08817_));
 sky130_fd_sc_hd__nor4_1 _16173_ (.A(_08816_),
    .B(_08075_),
    .C(_08817_),
    .D(_08784_),
    .Y(_08818_));
 sky130_fd_sc_hd__o22a_1 _16174_ (.A1(_08816_),
    .A2(_08075_),
    .B1(_08817_),
    .B2(_08784_),
    .X(_08819_));
 sky130_fd_sc_hd__or2_1 _16175_ (.A(_08818_),
    .B(_08819_),
    .X(_08820_));
 sky130_fd_sc_hd__clkbuf_4 _16176_ (.A(_08674_),
    .X(_08821_));
 sky130_fd_sc_hd__or3_1 _16177_ (.A(_08112_),
    .B(_08328_),
    .C(_08747_),
    .X(_08822_));
 sky130_fd_sc_hd__clkbuf_4 _16178_ (.A(_08112_),
    .X(_08823_));
 sky130_fd_sc_hd__o22ai_1 _16179_ (.A1(_08519_),
    .A2(_08823_),
    .B1(_08329_),
    .B2(_08377_),
    .Y(_08824_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(_08822_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__o31a_1 _16181_ (.A1(_08816_),
    .A2(_08821_),
    .A3(_08825_),
    .B1(_08822_),
    .X(_08826_));
 sky130_fd_sc_hd__xor2_1 _16182_ (.A(_08820_),
    .B(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__or2_1 _16183_ (.A(_08194_),
    .B(_08491_),
    .X(_08828_));
 sky130_fd_sc_hd__o22a_1 _16184_ (.A1(_08170_),
    .A2(_08042_),
    .B1(_08128_),
    .B2(_08180_),
    .X(_08829_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_07981_),
    .B(_08128_),
    .Y(_08830_));
 sky130_fd_sc_hd__nand2_1 _16186_ (.A(_08788_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__and2b_1 _16187_ (.A_N(_08829_),
    .B(_08831_),
    .X(_08832_));
 sky130_fd_sc_hd__xnor2_1 _16188_ (.A(_08828_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__nor2_1 _16189_ (.A(_08820_),
    .B(_08826_),
    .Y(_08834_));
 sky130_fd_sc_hd__a21oi_1 _16190_ (.A1(_08827_),
    .A2(_08833_),
    .B1(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__xor2_1 _16191_ (.A(_08815_),
    .B(_08835_),
    .X(_08836_));
 sky130_fd_sc_hd__or3b_1 _16192_ (.A(_08828_),
    .B(_08829_),
    .C_N(_08831_),
    .X(_08837_));
 sky130_fd_sc_hd__o21a_1 _16193_ (.A1(_08284_),
    .A2(_08579_),
    .B1(_08727_),
    .X(_08838_));
 sky130_fd_sc_hd__or2_1 _16194_ (.A(_08793_),
    .B(_08838_),
    .X(_08839_));
 sky130_fd_sc_hd__a21oi_1 _16195_ (.A1(_08831_),
    .A2(_08837_),
    .B1(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__and3_1 _16196_ (.A(_08831_),
    .B(_08837_),
    .C(_08839_),
    .X(_08841_));
 sky130_fd_sc_hd__nor2_1 _16197_ (.A(_08840_),
    .B(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__nor2_1 _16198_ (.A(_08815_),
    .B(_08835_),
    .Y(_08843_));
 sky130_fd_sc_hd__a21oi_1 _16199_ (.A1(_08836_),
    .A2(_08842_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__or2_1 _16200_ (.A(_08812_),
    .B(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__xor2_1 _16201_ (.A(_08812_),
    .B(_08844_),
    .X(_08846_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(_08840_),
    .B(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__and2b_1 _16203_ (.A_N(_08799_),
    .B(_08798_),
    .X(_08848_));
 sky130_fd_sc_hd__xnor2_1 _16204_ (.A(_08778_),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__a21o_1 _16205_ (.A1(_08845_),
    .A2(_08847_),
    .B1(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__inv_2 _16206_ (.A(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__or2_1 _16207_ (.A(_08840_),
    .B(_08846_),
    .X(_08852_));
 sky130_fd_sc_hd__nand2_1 _16208_ (.A(_08847_),
    .B(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__nor2_1 _16209_ (.A(_08519_),
    .B(_08053_),
    .Y(_08854_));
 sky130_fd_sc_hd__or3b_1 _16210_ (.A(_08377_),
    .B(_08329_),
    .C_N(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__nor2_1 _16211_ (.A(_08377_),
    .B(_08054_),
    .Y(_08856_));
 sky130_fd_sc_hd__a21o_1 _16212_ (.A1(_08227_),
    .A2(_08331_),
    .B1(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__nand2_1 _16213_ (.A(_08855_),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__nor2_1 _16214_ (.A(_08816_),
    .B(_08823_),
    .Y(_08859_));
 sky130_fd_sc_hd__xor2_1 _16215_ (.A(_08858_),
    .B(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__nor2_1 _16216_ (.A(_08377_),
    .B(_08062_),
    .Y(_08861_));
 sky130_fd_sc_hd__xor2_1 _16217_ (.A(_08854_),
    .B(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__and3_1 _16218_ (.A(_08250_),
    .B(_08331_),
    .C(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__a21oi_1 _16219_ (.A1(_08854_),
    .A2(_08861_),
    .B1(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__or2_1 _16220_ (.A(_08860_),
    .B(_08864_),
    .X(_08865_));
 sky130_fd_sc_hd__nand2_1 _16221_ (.A(_08860_),
    .B(_08864_),
    .Y(_08866_));
 sky130_fd_sc_hd__and2_1 _16222_ (.A(_08865_),
    .B(_08866_),
    .X(_08867_));
 sky130_fd_sc_hd__or2_1 _16223_ (.A(_08180_),
    .B(_08491_),
    .X(_08868_));
 sky130_fd_sc_hd__or2_1 _16224_ (.A(_08170_),
    .B(_08572_),
    .X(_08869_));
 sky130_fd_sc_hd__or2_1 _16225_ (.A(_08868_),
    .B(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__inv_2 _16226_ (.A(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__clkbuf_4 _16227_ (.A(_08170_),
    .X(_08872_));
 sky130_fd_sc_hd__clkbuf_4 _16228_ (.A(_08180_),
    .X(_08873_));
 sky130_fd_sc_hd__o22a_1 _16229_ (.A1(_08872_),
    .A2(_08491_),
    .B1(_08579_),
    .B2(_08873_),
    .X(_08874_));
 sky130_fd_sc_hd__nor2_1 _16230_ (.A(_08871_),
    .B(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__nand2_1 _16231_ (.A(_08867_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__or2_1 _16232_ (.A(_08194_),
    .B(_08579_),
    .X(_08877_));
 sky130_fd_sc_hd__xnor2_1 _16233_ (.A(_08830_),
    .B(_08868_),
    .Y(_08878_));
 sky130_fd_sc_hd__xnor2_1 _16234_ (.A(_08877_),
    .B(_08878_),
    .Y(_08879_));
 sky130_fd_sc_hd__nor2_1 _16235_ (.A(_08816_),
    .B(_08821_),
    .Y(_08880_));
 sky130_fd_sc_hd__xor2_1 _16236_ (.A(_08825_),
    .B(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__a21boi_1 _16237_ (.A1(_08857_),
    .A2(_08859_),
    .B1_N(_08855_),
    .Y(_08882_));
 sky130_fd_sc_hd__xor2_1 _16238_ (.A(_08881_),
    .B(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__xnor2_1 _16239_ (.A(_08879_),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__a21o_1 _16240_ (.A1(_08865_),
    .A2(_08876_),
    .B1(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__nand3_1 _16241_ (.A(_08884_),
    .B(_08865_),
    .C(_08876_),
    .Y(_08886_));
 sky130_fd_sc_hd__and2_1 _16242_ (.A(_08885_),
    .B(_08886_),
    .X(_08887_));
 sky130_fd_sc_hd__nand2_1 _16243_ (.A(_08871_),
    .B(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__xnor2_1 _16244_ (.A(_08827_),
    .B(_08833_),
    .Y(_08889_));
 sky130_fd_sc_hd__nor2_1 _16245_ (.A(_08881_),
    .B(_08882_),
    .Y(_08890_));
 sky130_fd_sc_hd__a21oi_1 _16246_ (.A1(_08879_),
    .A2(_08883_),
    .B1(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__xor2_1 _16247_ (.A(_08889_),
    .B(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__or3_1 _16248_ (.A(_08872_),
    .B(_08128_),
    .C(_08868_),
    .X(_08893_));
 sky130_fd_sc_hd__or2b_1 _16249_ (.A(_08877_),
    .B_N(_08878_),
    .X(_08894_));
 sky130_fd_sc_hd__clkbuf_4 _16250_ (.A(_08283_),
    .X(_08895_));
 sky130_fd_sc_hd__or2_1 _16251_ (.A(_08895_),
    .B(_08579_),
    .X(_08896_));
 sky130_fd_sc_hd__a21oi_1 _16252_ (.A1(_08893_),
    .A2(_08894_),
    .B1(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__and3_1 _16253_ (.A(_08896_),
    .B(_08893_),
    .C(_08894_),
    .X(_08898_));
 sky130_fd_sc_hd__nor2_1 _16254_ (.A(_08897_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__xnor2_1 _16255_ (.A(_08892_),
    .B(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__a21oi_1 _16256_ (.A1(_08885_),
    .A2(_08888_),
    .B1(_08900_),
    .Y(_08901_));
 sky130_fd_sc_hd__xnor2_1 _16257_ (.A(_08836_),
    .B(_08842_),
    .Y(_08902_));
 sky130_fd_sc_hd__nor2_1 _16258_ (.A(_08889_),
    .B(_08891_),
    .Y(_08903_));
 sky130_fd_sc_hd__a21oi_1 _16259_ (.A1(_08892_),
    .A2(_08899_),
    .B1(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__nor2_1 _16260_ (.A(_08902_),
    .B(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(_08902_),
    .B(_08904_),
    .Y(_08906_));
 sky130_fd_sc_hd__and2b_1 _16262_ (.A_N(_08905_),
    .B(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__xor2_1 _16263_ (.A(_08897_),
    .B(_08907_),
    .X(_08908_));
 sky130_fd_sc_hd__a21o_1 _16264_ (.A1(_08897_),
    .A2(_08906_),
    .B1(_08905_),
    .X(_08909_));
 sky130_fd_sc_hd__a21oi_1 _16265_ (.A1(_08901_),
    .A2(_08908_),
    .B1(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__nor2_1 _16266_ (.A(_08853_),
    .B(_08910_),
    .Y(_08911_));
 sky130_fd_sc_hd__or4_1 _16267_ (.A(_08226_),
    .B(_08816_),
    .C(_08162_),
    .D(_08160_),
    .X(_08912_));
 sky130_fd_sc_hd__a21o_1 _16268_ (.A1(_08215_),
    .A2(_08335_),
    .B1(_08856_),
    .X(_08913_));
 sky130_fd_sc_hd__a21oi_1 _16269_ (.A1(_08250_),
    .A2(_08331_),
    .B1(_08862_),
    .Y(_08914_));
 sky130_fd_sc_hd__or2_1 _16270_ (.A(_08863_),
    .B(_08914_),
    .X(_08915_));
 sky130_fd_sc_hd__o22a_1 _16271_ (.A1(_08215_),
    .A2(_08162_),
    .B1(_08160_),
    .B2(_08226_),
    .X(_08916_));
 sky130_fd_sc_hd__or4_1 _16272_ (.A(_08215_),
    .B(_08226_),
    .C(_08135_),
    .D(_08160_),
    .X(_08917_));
 sky130_fd_sc_hd__o31ai_2 _16273_ (.A1(_08816_),
    .A2(_08335_),
    .A3(_08916_),
    .B1(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__xor2_1 _16274_ (.A(_08915_),
    .B(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__nand2_1 _16275_ (.A(_08869_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__or2_1 _16276_ (.A(_08869_),
    .B(_08919_),
    .X(_08921_));
 sky130_fd_sc_hd__and4b_1 _16277_ (.A_N(_08912_),
    .B(_08913_),
    .C(_08920_),
    .D(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__or2_1 _16278_ (.A(_08867_),
    .B(_08875_),
    .X(_08923_));
 sky130_fd_sc_hd__nand2_1 _16279_ (.A(_08876_),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__inv_2 _16280_ (.A(_08918_),
    .Y(_08925_));
 sky130_fd_sc_hd__o21a_1 _16281_ (.A1(_08915_),
    .A2(_08925_),
    .B1(_08921_),
    .X(_08926_));
 sky130_fd_sc_hd__nor2_1 _16282_ (.A(_08924_),
    .B(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__nand2_1 _16283_ (.A(_08924_),
    .B(_08926_),
    .Y(_08928_));
 sky130_fd_sc_hd__xnor2_1 _16284_ (.A(_08870_),
    .B(_08887_),
    .Y(_08929_));
 sky130_fd_sc_hd__o211a_1 _16285_ (.A1(_08922_),
    .A2(_08927_),
    .B1(_08928_),
    .C1(_08929_),
    .X(_08930_));
 sky130_fd_sc_hd__or2b_1 _16286_ (.A(_08909_),
    .B_N(_08853_),
    .X(_08931_));
 sky130_fd_sc_hd__and3_1 _16287_ (.A(_08900_),
    .B(_08885_),
    .C(_08888_),
    .X(_08932_));
 sky130_fd_sc_hd__nor2_1 _16288_ (.A(_08901_),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__and4_1 _16289_ (.A(_08908_),
    .B(_08930_),
    .C(_08931_),
    .D(_08933_),
    .X(_08934_));
 sky130_fd_sc_hd__and3_1 _16290_ (.A(_08849_),
    .B(_08845_),
    .C(_08847_),
    .X(_08935_));
 sky130_fd_sc_hd__o21ba_1 _16291_ (.A1(_08911_),
    .A2(_08934_),
    .B1_N(_08935_),
    .X(_08936_));
 sky130_fd_sc_hd__xor2_1 _16292_ (.A(_08764_),
    .B(_08807_),
    .X(_08937_));
 sky130_fd_sc_hd__a21bo_1 _16293_ (.A1(_08806_),
    .A2(_08801_),
    .B1_N(_08805_),
    .X(_08938_));
 sky130_fd_sc_hd__a211oi_1 _16294_ (.A1(_08803_),
    .A2(_08804_),
    .B1(_08807_),
    .C1(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__o211a_1 _16295_ (.A1(_08851_),
    .A2(_08936_),
    .B1(_08937_),
    .C1(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__nor2_1 _16296_ (.A(_08719_),
    .B(_08763_),
    .Y(_08941_));
 sky130_fd_sc_hd__a21oi_1 _16297_ (.A1(_08764_),
    .A2(_08807_),
    .B1(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__xnor2_2 _16298_ (.A(_08811_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__a32oi_4 _16299_ (.A1(_08764_),
    .A2(_08807_),
    .A3(_08811_),
    .B1(_08940_),
    .B2(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__xnor2_1 _16300_ (.A(_08620_),
    .B(_08670_),
    .Y(_08945_));
 sky130_fd_sc_hd__nor2_1 _16301_ (.A(_08808_),
    .B(_08810_),
    .Y(_08946_));
 sky130_fd_sc_hd__a21oi_1 _16302_ (.A1(_08941_),
    .A2(_08811_),
    .B1(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__xnor2_1 _16303_ (.A(_08945_),
    .B(_08947_),
    .Y(_08948_));
 sky130_fd_sc_hd__and2_1 _16304_ (.A(_08941_),
    .B(_08811_),
    .X(_08949_));
 sky130_fd_sc_hd__inv_2 _16305_ (.A(_08945_),
    .Y(_08950_));
 sky130_fd_sc_hd__a2bb2o_2 _16306_ (.A1_N(_08944_),
    .A2_N(_08948_),
    .B1(_08949_),
    .B2(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__a21o_1 _16307_ (.A1(_08950_),
    .A2(_08946_),
    .B1(_08671_),
    .X(_08952_));
 sky130_fd_sc_hd__xnor2_4 _16308_ (.A(_08619_),
    .B(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__and3b_1 _16309_ (.A_N(_08619_),
    .B(_08950_),
    .C(_08946_),
    .X(_08954_));
 sky130_fd_sc_hd__a21oi_4 _16310_ (.A1(_08951_),
    .A2(_08953_),
    .B1(_08954_),
    .Y(_08955_));
 sky130_fd_sc_hd__nand2_1 _16311_ (.A(_08617_),
    .B(_08672_),
    .Y(_08956_));
 sky130_fd_sc_hd__o221ai_4 _16312_ (.A1(_08550_),
    .A2(_08616_),
    .B1(_08673_),
    .B2(_08955_),
    .C1(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__or3_1 _16313_ (.A(_08292_),
    .B(_07996_),
    .C(_07959_),
    .X(_08958_));
 sky130_fd_sc_hd__a21bo_1 _16314_ (.A1(_08290_),
    .A2(_08291_),
    .B1_N(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__or2_1 _16315_ (.A(_08008_),
    .B(_08204_),
    .X(_08960_));
 sky130_fd_sc_hd__a2bb2o_1 _16316_ (.A1_N(_08192_),
    .A2_N(_08960_),
    .B1(_08179_),
    .B2(_08190_),
    .X(_08961_));
 sky130_fd_sc_hd__nor2_1 _16317_ (.A(_07924_),
    .B(_08276_),
    .Y(_08962_));
 sky130_fd_sc_hd__and2b_1 _16318_ (.A_N(_07913_),
    .B(_08264_),
    .X(_08963_));
 sky130_fd_sc_hd__xnor2_1 _16319_ (.A(_08962_),
    .B(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__nor2_1 _16320_ (.A(_08282_),
    .B(_07959_),
    .Y(_08965_));
 sky130_fd_sc_hd__xnor2_1 _16321_ (.A(_08964_),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__xor2_1 _16322_ (.A(_08961_),
    .B(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__nand2_1 _16323_ (.A(_08959_),
    .B(_08967_),
    .Y(_08968_));
 sky130_fd_sc_hd__or2_1 _16324_ (.A(_08959_),
    .B(_08967_),
    .X(_08969_));
 sky130_fd_sc_hd__and2_2 _16325_ (.A(_08968_),
    .B(_08969_),
    .X(_08970_));
 sky130_fd_sc_hd__a21boi_2 _16326_ (.A1(_05209_),
    .A2(\rbzero.wall_tracer.stepDistX[3] ),
    .B1_N(_08214_),
    .Y(_08971_));
 sky130_fd_sc_hd__o22a_1 _16327_ (.A1(_08180_),
    .A2(_08189_),
    .B1(_08971_),
    .B2(_08170_),
    .X(_08972_));
 sky130_fd_sc_hd__or4_1 _16328_ (.A(_07981_),
    .B(_07989_),
    .C(_08189_),
    .D(_08971_),
    .X(_08973_));
 sky130_fd_sc_hd__or2b_1 _16329_ (.A(_08972_),
    .B_N(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__nor2_1 _16330_ (.A(_08178_),
    .B(_08194_),
    .Y(_08975_));
 sky130_fd_sc_hd__xnor2_2 _16331_ (.A(_08974_),
    .B(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__or4b_2 _16332_ (.A(_07602_),
    .B(_08230_),
    .C(_08147_),
    .D_N(_08225_),
    .X(_08977_));
 sky130_fd_sc_hd__or4_1 _16333_ (.A(_07598_),
    .B(_08230_),
    .C(_08147_),
    .D(_08236_),
    .X(_08978_));
 sky130_fd_sc_hd__xnor2_2 _16334_ (.A(_08977_),
    .B(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__nand2_1 _16335_ (.A(_08230_),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_08980_));
 sky130_fd_sc_hd__inv_2 _16336_ (.A(_07571_),
    .Y(_08981_));
 sky130_fd_sc_hd__a31o_1 _16337_ (.A1(_08218_),
    .A2(_08232_),
    .A3(_08208_),
    .B1(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__or4_2 _16338_ (.A(_07566_),
    .B(_07568_),
    .C(_07571_),
    .D(_08220_),
    .X(_08983_));
 sky130_fd_sc_hd__a31o_1 _16339_ (.A1(_05194_),
    .A2(_08982_),
    .A3(_08983_),
    .B1(_08224_),
    .X(_08984_));
 sky130_fd_sc_hd__a21o_1 _16340_ (.A1(_08980_),
    .A2(_08984_),
    .B1(_08147_),
    .X(_08985_));
 sky130_fd_sc_hd__nor2_1 _16341_ (.A(_08239_),
    .B(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__xnor2_2 _16342_ (.A(_08979_),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__or2_1 _16343_ (.A(_08977_),
    .B(_08243_),
    .X(_08988_));
 sky130_fd_sc_hd__o31a_1 _16344_ (.A1(_08237_),
    .A2(_08239_),
    .A3(_08229_),
    .B1(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__xnor2_2 _16345_ (.A(_08987_),
    .B(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__xnor2_2 _16346_ (.A(_08976_),
    .B(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__nor2_1 _16347_ (.A(_08241_),
    .B(_08247_),
    .Y(_08992_));
 sky130_fd_sc_hd__a21o_1 _16348_ (.A1(_08206_),
    .A2(_08248_),
    .B1(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__xnor2_2 _16349_ (.A(_08991_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__xnor2_4 _16350_ (.A(_08970_),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(_08249_),
    .B(_08280_),
    .Y(_08996_));
 sky130_fd_sc_hd__a21oi_4 _16352_ (.A1(_08281_),
    .A2(_08296_),
    .B1(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__xor2_4 _16353_ (.A(_08995_),
    .B(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__nor2_1 _16354_ (.A(_08363_),
    .B(_08364_),
    .Y(_08999_));
 sky130_fd_sc_hd__a21o_2 _16355_ (.A1(_08358_),
    .A2(_08365_),
    .B1(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__or2b_1 _16356_ (.A(_08295_),
    .B_N(_08288_),
    .X(_09001_));
 sky130_fd_sc_hd__a21bo_1 _16357_ (.A1(_08289_),
    .A2(_08294_),
    .B1_N(_09001_),
    .X(_09002_));
 sky130_fd_sc_hd__or4_1 _16358_ (.A(_07967_),
    .B(_08674_),
    .C(_08034_),
    .D(_08045_),
    .X(_09003_));
 sky130_fd_sc_hd__o22ai_1 _16359_ (.A1(_07967_),
    .A2(_08035_),
    .B1(_08046_),
    .B2(_08674_),
    .Y(_09004_));
 sky130_fd_sc_hd__nand2_1 _16360_ (.A(_09003_),
    .B(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__or3_1 _16361_ (.A(_08823_),
    .B(_08058_),
    .C(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__o21ai_1 _16362_ (.A1(_08823_),
    .A2(_08059_),
    .B1(_09005_),
    .Y(_09007_));
 sky130_fd_sc_hd__and2_1 _16363_ (.A(_09006_),
    .B(_09007_),
    .X(_09008_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_07995_),
    .B(_08570_),
    .Y(_09009_));
 sky130_fd_sc_hd__o22a_1 _16365_ (.A1(_07995_),
    .A2(_08109_),
    .B1(_08084_),
    .B2(_07931_),
    .X(_09010_));
 sky130_fd_sc_hd__a21o_1 _16366_ (.A1(_08360_),
    .A2(_09009_),
    .B1(_09010_),
    .X(_09011_));
 sky130_fd_sc_hd__or2_1 _16367_ (.A(_07941_),
    .B(_08097_),
    .X(_09012_));
 sky130_fd_sc_hd__xnor2_1 _16368_ (.A(_09011_),
    .B(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__nand2_1 _16369_ (.A(_08359_),
    .B(_08360_),
    .Y(_09014_));
 sky130_fd_sc_hd__o31a_1 _16370_ (.A1(_08361_),
    .A2(_07967_),
    .A3(_08097_),
    .B1(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__nor2_1 _16371_ (.A(_09013_),
    .B(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__and2_1 _16372_ (.A(_09013_),
    .B(_09015_),
    .X(_09017_));
 sky130_fd_sc_hd__nor2_1 _16373_ (.A(_09016_),
    .B(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__xor2_2 _16374_ (.A(_09008_),
    .B(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__xnor2_2 _16375_ (.A(_09002_),
    .B(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__xnor2_4 _16376_ (.A(_09000_),
    .B(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__xnor2_4 _16377_ (.A(_08998_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__nor2_1 _16378_ (.A(_08297_),
    .B(_08326_),
    .Y(_09023_));
 sky130_fd_sc_hd__a21oi_4 _16379_ (.A1(_08327_),
    .A2(_08370_),
    .B1(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__xor2_4 _16380_ (.A(_09022_),
    .B(_09024_),
    .X(_09025_));
 sky130_fd_sc_hd__or2b_1 _16381_ (.A(_08369_),
    .B_N(_08349_),
    .X(_09026_));
 sky130_fd_sc_hd__nand2_8 _16382_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08148_),
    .Y(_09027_));
 sky130_fd_sc_hd__or2_2 _16383_ (.A(_08147_),
    .B(_09027_),
    .X(_09028_));
 sky130_fd_sc_hd__clkbuf_4 _16384_ (.A(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__nor2_2 _16385_ (.A(_09029_),
    .B(_08162_),
    .Y(_09030_));
 sky130_fd_sc_hd__a21bo_1 _16386_ (.A1(_08416_),
    .A2(_08420_),
    .B1_N(_08426_),
    .X(_09031_));
 sky130_fd_sc_hd__nand2_1 _16387_ (.A(_08331_),
    .B(_08420_),
    .Y(_09032_));
 sky130_fd_sc_hd__a2bb2o_1 _16388_ (.A1_N(_08053_),
    .A2_N(_08158_),
    .B1(_08418_),
    .B2(_08039_),
    .X(_09033_));
 sky130_fd_sc_hd__nand2_1 _16389_ (.A(_09032_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__nor2_1 _16390_ (.A(_08062_),
    .B(_08425_),
    .Y(_09035_));
 sky130_fd_sc_hd__xor2_1 _16391_ (.A(_09034_),
    .B(_09035_),
    .X(_09036_));
 sky130_fd_sc_hd__a21oi_1 _16392_ (.A1(_08352_),
    .A2(_08355_),
    .B1(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__and3_1 _16393_ (.A(_08352_),
    .B(_08355_),
    .C(_09036_),
    .X(_09038_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(_09037_),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__xnor2_2 _16395_ (.A(_09031_),
    .B(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__nor2_1 _16396_ (.A(_08161_),
    .B(_08431_),
    .Y(_09041_));
 sky130_fd_sc_hd__nor2_1 _16397_ (.A(_08430_),
    .B(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__xnor2_1 _16398_ (.A(_09040_),
    .B(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__xnor2_1 _16399_ (.A(_09030_),
    .B(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__a21o_1 _16400_ (.A1(_08367_),
    .A2(_09026_),
    .B1(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__nand3_2 _16401_ (.A(_08367_),
    .B(_09026_),
    .C(_09044_),
    .Y(_09046_));
 sky130_fd_sc_hd__nand2_2 _16402_ (.A(_09045_),
    .B(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__and2_2 _16403_ (.A(_08165_),
    .B(_08432_),
    .X(_09048_));
 sky130_fd_sc_hd__xnor2_4 _16404_ (.A(_09047_),
    .B(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__xnor2_4 _16405_ (.A(_09025_),
    .B(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__nor2_1 _16406_ (.A(_08371_),
    .B(_08411_),
    .Y(_09051_));
 sky130_fd_sc_hd__a21oi_2 _16407_ (.A1(_08412_),
    .A2(_08438_),
    .B1(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__xor2_2 _16408_ (.A(_09050_),
    .B(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__inv_2 _16409_ (.A(_08437_),
    .Y(_09054_));
 sky130_fd_sc_hd__o21a_1 _16410_ (.A1(_08413_),
    .A2(_09054_),
    .B1(_08435_),
    .X(_09055_));
 sky130_fd_sc_hd__xnor2_2 _16411_ (.A(_09053_),
    .B(_09055_),
    .Y(_09056_));
 sky130_fd_sc_hd__nor2_1 _16412_ (.A(_08439_),
    .B(_08468_),
    .Y(_09057_));
 sky130_fd_sc_hd__a21o_1 _16413_ (.A1(_08169_),
    .A2(_08469_),
    .B1(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__xnor2_2 _16414_ (.A(_09056_),
    .B(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__xnor2_2 _16415_ (.A(_09059_),
    .B(_08547_),
    .Y(_09060_));
 sky130_fd_sc_hd__a21o_2 _16416_ (.A1(_08549_),
    .A2(_08957_),
    .B1(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__nand3_4 _16417_ (.A(_08549_),
    .B(_08957_),
    .C(_09060_),
    .Y(_09062_));
 sky130_fd_sc_hd__mux2_1 _16418_ (.A0(\rbzero.debug_overlay.playerY[-6] ),
    .A1(\rbzero.debug_overlay.playerX[-6] ),
    .S(_07895_),
    .X(_09063_));
 sky130_fd_sc_hd__and3_1 _16419_ (.A(_09061_),
    .B(_09062_),
    .C(_09063_),
    .X(_09064_));
 sky130_fd_sc_hd__a21o_1 _16420_ (.A1(_09061_),
    .A2(_09062_),
    .B1(_09063_),
    .X(_09065_));
 sky130_fd_sc_hd__or2b_1 _16421_ (.A(_09064_),
    .B_N(_09065_),
    .X(_09066_));
 sky130_fd_sc_hd__xor2_2 _16422_ (.A(_08617_),
    .B(_08672_),
    .X(_09067_));
 sky130_fd_sc_hd__xnor2_4 _16423_ (.A(_09067_),
    .B(_08955_),
    .Y(_09068_));
 sky130_fd_sc_hd__xor2_4 _16424_ (.A(_08951_),
    .B(_08953_),
    .X(_09069_));
 sky130_fd_sc_hd__mux2_1 _16425_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_07894_),
    .X(_09070_));
 sky130_fd_sc_hd__mux2_1 _16426_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_07895_),
    .X(_09071_));
 sky130_fd_sc_hd__a21o_1 _16427_ (.A1(_09069_),
    .A2(_09070_),
    .B1(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__and3_1 _16428_ (.A(_09071_),
    .B(_09069_),
    .C(_09070_),
    .X(_09073_));
 sky130_fd_sc_hd__a21o_1 _16429_ (.A1(_09068_),
    .A2(_09072_),
    .B1(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__mux2_1 _16430_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_07895_),
    .X(_09075_));
 sky130_fd_sc_hd__xor2_4 _16431_ (.A(_08549_),
    .B(_08957_),
    .X(_09076_));
 sky130_fd_sc_hd__a21o_1 _16432_ (.A1(_09074_),
    .A2(_09075_),
    .B1(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__or2_1 _16433_ (.A(_09074_),
    .B(_09075_),
    .X(_09078_));
 sky130_fd_sc_hd__nand2_1 _16434_ (.A(_09077_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__xor2_2 _16435_ (.A(_09066_),
    .B(_09079_),
    .X(_09080_));
 sky130_fd_sc_hd__mux2_1 _16436_ (.A0(_05397_),
    .A1(_05503_),
    .S(_07971_),
    .X(_09081_));
 sky130_fd_sc_hd__buf_4 _16437_ (.A(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__nor2_1 _16438_ (.A(_09080_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__a21o_1 _16439_ (.A1(_09080_),
    .A2(_09082_),
    .B1(_05194_),
    .X(_09084_));
 sky130_fd_sc_hd__buf_4 _16440_ (.A(_07970_),
    .X(_09085_));
 sky130_fd_sc_hd__or2_1 _16441_ (.A(\rbzero.wall_tracer.texu[0] ),
    .B(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__o211a_1 _16442_ (.A1(_09083_),
    .A2(_09084_),
    .B1(_09086_),
    .C1(_07642_),
    .X(_00511_));
 sky130_fd_sc_hd__and2b_1 _16443_ (.A_N(_09059_),
    .B(_08547_),
    .X(_09087_));
 sky130_fd_sc_hd__a31o_1 _16444_ (.A1(_08549_),
    .A2(_08957_),
    .A3(_09060_),
    .B1(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__nand2_1 _16445_ (.A(_09056_),
    .B(_09058_),
    .Y(_09089_));
 sky130_fd_sc_hd__a21o_1 _16446_ (.A1(_09008_),
    .A2(_09018_),
    .B1(_09016_),
    .X(_09090_));
 sky130_fd_sc_hd__nand2_1 _16447_ (.A(_08961_),
    .B(_08966_),
    .Y(_09091_));
 sky130_fd_sc_hd__or4_1 _16448_ (.A(_07941_),
    .B(_08075_),
    .C(_08035_),
    .D(_08046_),
    .X(_09092_));
 sky130_fd_sc_hd__o22ai_1 _16449_ (.A1(_07941_),
    .A2(_08035_),
    .B1(_08046_),
    .B2(_08075_),
    .Y(_09093_));
 sky130_fd_sc_hd__nand2_1 _16450_ (.A(_09092_),
    .B(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__or3_1 _16451_ (.A(_08821_),
    .B(_08059_),
    .C(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__clkbuf_4 _16452_ (.A(_08821_),
    .X(_09096_));
 sky130_fd_sc_hd__o21ai_1 _16453_ (.A1(_09096_),
    .A2(_08356_),
    .B1(_09094_),
    .Y(_09097_));
 sky130_fd_sc_hd__and2_1 _16454_ (.A(_09095_),
    .B(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__nor2_1 _16455_ (.A(_07977_),
    .B(_08109_),
    .Y(_09099_));
 sky130_fd_sc_hd__xnor2_1 _16456_ (.A(_09009_),
    .B(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__or2_1 _16457_ (.A(_07932_),
    .B(_08097_),
    .X(_09101_));
 sky130_fd_sc_hd__xnor2_1 _16458_ (.A(_09100_),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__clkbuf_4 _16459_ (.A(_08097_),
    .X(_09103_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(_08360_),
    .B(_09009_),
    .Y(_09104_));
 sky130_fd_sc_hd__o31a_1 _16461_ (.A1(_07941_),
    .A2(_09103_),
    .A3(_09010_),
    .B1(_09104_),
    .X(_09105_));
 sky130_fd_sc_hd__nor2_1 _16462_ (.A(_09102_),
    .B(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__and2_1 _16463_ (.A(_09102_),
    .B(_09105_),
    .X(_09107_));
 sky130_fd_sc_hd__nor2_1 _16464_ (.A(_09106_),
    .B(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__xnor2_1 _16465_ (.A(_09098_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__a21oi_1 _16466_ (.A1(_09091_),
    .A2(_08968_),
    .B1(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__and3_1 _16467_ (.A(_09091_),
    .B(_08968_),
    .C(_09109_),
    .X(_09111_));
 sky130_fd_sc_hd__nor2_1 _16468_ (.A(_09110_),
    .B(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__xor2_2 _16469_ (.A(_09090_),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__clkbuf_4 _16470_ (.A(_07959_),
    .X(_09114_));
 sky130_fd_sc_hd__or3_1 _16471_ (.A(_08282_),
    .B(_09114_),
    .C(_08964_),
    .X(_09115_));
 sky130_fd_sc_hd__a21bo_1 _16472_ (.A1(_08962_),
    .A2(_08963_),
    .B1_N(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__buf_4 _16473_ (.A(_08194_),
    .X(_09117_));
 sky130_fd_sc_hd__o31ai_2 _16474_ (.A1(_08178_),
    .A2(_09117_),
    .A3(_08972_),
    .B1(_08973_),
    .Y(_09118_));
 sky130_fd_sc_hd__nor2_2 _16475_ (.A(_08284_),
    .B(_08177_),
    .Y(_09119_));
 sky130_fd_sc_hd__a2bb2o_1 _16476_ (.A1_N(_08283_),
    .A2_N(_08177_),
    .B1(_08264_),
    .B2(_08626_),
    .X(_09120_));
 sky130_fd_sc_hd__a21bo_1 _16477_ (.A1(_08963_),
    .A2(_09119_),
    .B1_N(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__nor2_1 _16478_ (.A(_08383_),
    .B(_07959_),
    .Y(_09122_));
 sky130_fd_sc_hd__xnor2_1 _16479_ (.A(_09121_),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__xnor2_1 _16480_ (.A(_09118_),
    .B(_09123_),
    .Y(_09124_));
 sky130_fd_sc_hd__xnor2_2 _16481_ (.A(_09116_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__clkbuf_4 _16482_ (.A(_08189_),
    .X(_09126_));
 sky130_fd_sc_hd__nor2_1 _16483_ (.A(_09126_),
    .B(_08194_),
    .Y(_09127_));
 sky130_fd_sc_hd__nor2_1 _16484_ (.A(_08180_),
    .B(_08971_),
    .Y(_09128_));
 sky130_fd_sc_hd__nand2_2 _16485_ (.A(_05209_),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_09129_));
 sky130_fd_sc_hd__a21oi_2 _16486_ (.A1(_08242_),
    .A2(_09129_),
    .B1(_08170_),
    .Y(_09130_));
 sky130_fd_sc_hd__xor2_2 _16487_ (.A(_09128_),
    .B(_09130_),
    .X(_09131_));
 sky130_fd_sc_hd__xor2_2 _16488_ (.A(_09127_),
    .B(_09131_),
    .X(_09132_));
 sky130_fd_sc_hd__or4_1 _16489_ (.A(_07602_),
    .B(_08230_),
    .C(_08147_),
    .D(_08236_),
    .X(_09133_));
 sky130_fd_sc_hd__or4_1 _16490_ (.A(_07598_),
    .B(_08230_),
    .C(_08147_),
    .D(_08984_),
    .X(_09134_));
 sky130_fd_sc_hd__xnor2_1 _16491_ (.A(_09133_),
    .B(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__o41a_1 _16492_ (.A1(_07566_),
    .A2(_07568_),
    .A3(_07571_),
    .A4(_08220_),
    .B1(_07575_),
    .X(_09136_));
 sky130_fd_sc_hd__a311o_1 _16493_ (.A1(_08981_),
    .A2(_07574_),
    .A3(_08234_),
    .B1(_09136_),
    .C1(_07970_),
    .X(_09137_));
 sky130_fd_sc_hd__a22oi_4 _16494_ (.A1(_08230_),
    .A2(\rbzero.wall_tracer.stepDistY[7] ),
    .B1(_08235_),
    .B2(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__nor2_1 _16495_ (.A(_08816_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__xnor2_1 _16496_ (.A(_09135_),
    .B(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__clkbuf_4 _16497_ (.A(_08985_),
    .X(_09141_));
 sky130_fd_sc_hd__or2_1 _16498_ (.A(_08977_),
    .B(_08978_),
    .X(_09142_));
 sky130_fd_sc_hd__o31a_1 _16499_ (.A1(_08979_),
    .A2(_08239_),
    .A3(_09141_),
    .B1(_09142_),
    .X(_09143_));
 sky130_fd_sc_hd__xnor2_2 _16500_ (.A(_09140_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__xnor2_2 _16501_ (.A(_09132_),
    .B(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__and2b_1 _16502_ (.A_N(_08989_),
    .B(_08987_),
    .X(_09146_));
 sky130_fd_sc_hd__a21oi_2 _16503_ (.A1(_08976_),
    .A2(_08990_),
    .B1(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__xor2_2 _16504_ (.A(_09145_),
    .B(_09147_),
    .X(_09148_));
 sky130_fd_sc_hd__xnor2_2 _16505_ (.A(_09125_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__or2b_1 _16506_ (.A(_08991_),
    .B_N(_08993_),
    .X(_09150_));
 sky130_fd_sc_hd__a21bo_1 _16507_ (.A1(_08970_),
    .A2(_08994_),
    .B1_N(_09150_),
    .X(_09151_));
 sky130_fd_sc_hd__xnor2_2 _16508_ (.A(_09149_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__xnor2_2 _16509_ (.A(_09113_),
    .B(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__nor2_1 _16510_ (.A(_08995_),
    .B(_08997_),
    .Y(_09154_));
 sky130_fd_sc_hd__a21oi_2 _16511_ (.A1(_08998_),
    .A2(_09021_),
    .B1(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__xor2_2 _16512_ (.A(_09153_),
    .B(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__nand2_1 _16513_ (.A(_09030_),
    .B(_09043_),
    .Y(_09157_));
 sky130_fd_sc_hd__o31ai_4 _16514_ (.A1(_09040_),
    .A2(_08430_),
    .A3(_09041_),
    .B1(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__or2b_1 _16515_ (.A(_09020_),
    .B_N(_09000_),
    .X(_09159_));
 sky130_fd_sc_hd__a21bo_1 _16516_ (.A1(_09002_),
    .A2(_09019_),
    .B1_N(_09159_),
    .X(_09160_));
 sky130_fd_sc_hd__and4_1 _16517_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_04015_),
    .C(_09030_),
    .D(_08416_),
    .X(_09161_));
 sky130_fd_sc_hd__nand2_4 _16518_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_04015_),
    .Y(_09162_));
 sky130_fd_sc_hd__or2_1 _16519_ (.A(_05209_),
    .B(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__buf_2 _16520_ (.A(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__clkbuf_4 _16521_ (.A(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__o22a_1 _16522_ (.A1(_09029_),
    .A2(_08160_),
    .B1(_09165_),
    .B2(_08162_),
    .X(_09166_));
 sky130_fd_sc_hd__a21bo_1 _16523_ (.A1(_09033_),
    .A2(_09035_),
    .B1_N(_09032_),
    .X(_09167_));
 sky130_fd_sc_hd__nand2_1 _16524_ (.A(_09003_),
    .B(_09006_),
    .Y(_09168_));
 sky130_fd_sc_hd__or3_1 _16525_ (.A(_08112_),
    .B(_08329_),
    .C(_08419_),
    .X(_09169_));
 sky130_fd_sc_hd__a2bb2o_1 _16526_ (.A1_N(_08112_),
    .A2_N(_08150_),
    .B1(_08331_),
    .B2(_08417_),
    .X(_09170_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(_09169_),
    .B(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__nor2_1 _16528_ (.A(_08054_),
    .B(_08425_),
    .Y(_09172_));
 sky130_fd_sc_hd__xor2_1 _16529_ (.A(_09171_),
    .B(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__xnor2_1 _16530_ (.A(_09168_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__xnor2_1 _16531_ (.A(_09167_),
    .B(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__a21oi_2 _16532_ (.A1(_09031_),
    .A2(_09039_),
    .B1(_09037_),
    .Y(_09176_));
 sky130_fd_sc_hd__xor2_1 _16533_ (.A(_09175_),
    .B(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__or3b_1 _16534_ (.A(_09161_),
    .B(_09166_),
    .C_N(_09177_),
    .X(_09178_));
 sky130_fd_sc_hd__o21bai_1 _16535_ (.A1(_09161_),
    .A2(_09166_),
    .B1_N(_09177_),
    .Y(_09179_));
 sky130_fd_sc_hd__and2_1 _16536_ (.A(_09178_),
    .B(_09179_),
    .X(_09180_));
 sky130_fd_sc_hd__xnor2_1 _16537_ (.A(_09160_),
    .B(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__xnor2_2 _16538_ (.A(_09158_),
    .B(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__xnor2_2 _16539_ (.A(_09156_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__nor2_1 _16540_ (.A(_09022_),
    .B(_09024_),
    .Y(_09184_));
 sky130_fd_sc_hd__a21oi_4 _16541_ (.A1(_09025_),
    .A2(_09049_),
    .B1(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__xnor2_4 _16542_ (.A(_09183_),
    .B(_09185_),
    .Y(_09186_));
 sky130_fd_sc_hd__a21boi_4 _16543_ (.A1(_09046_),
    .A2(_09048_),
    .B1_N(_09045_),
    .Y(_09187_));
 sky130_fd_sc_hd__xnor2_4 _16544_ (.A(_09186_),
    .B(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__inv_2 _16545_ (.A(_09055_),
    .Y(_09189_));
 sky130_fd_sc_hd__nor2_1 _16546_ (.A(_09050_),
    .B(_09052_),
    .Y(_09190_));
 sky130_fd_sc_hd__a21oi_2 _16547_ (.A1(_09053_),
    .A2(_09189_),
    .B1(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__xor2_2 _16548_ (.A(_09188_),
    .B(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__xnor2_2 _16549_ (.A(_09089_),
    .B(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__xnor2_4 _16550_ (.A(_09088_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__or2_1 _16551_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_07895_),
    .X(_09195_));
 sky130_fd_sc_hd__o21ai_2 _16552_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_07971_),
    .B1(_09195_),
    .Y(_09196_));
 sky130_fd_sc_hd__nor2_1 _16553_ (.A(_09194_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__nand2_1 _16554_ (.A(_09194_),
    .B(_09196_),
    .Y(_09198_));
 sky130_fd_sc_hd__or2b_1 _16555_ (.A(_09197_),
    .B_N(_09198_),
    .X(_09199_));
 sky130_fd_sc_hd__a31o_1 _16556_ (.A1(_09065_),
    .A2(_09077_),
    .A3(_09078_),
    .B1(_09064_),
    .X(_09200_));
 sky130_fd_sc_hd__xnor2_1 _16557_ (.A(_09199_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__xnor2_1 _16558_ (.A(_09082_),
    .B(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__or2_1 _16559_ (.A(\rbzero.wall_tracer.texu[1] ),
    .B(_09085_),
    .X(_09203_));
 sky130_fd_sc_hd__o211a_1 _16560_ (.A1(_05194_),
    .A2(_09202_),
    .B1(_09203_),
    .C1(_07642_),
    .X(_00512_));
 sky130_fd_sc_hd__and2b_1 _16561_ (.A_N(_09059_),
    .B(_09193_),
    .X(_09204_));
 sky130_fd_sc_hd__or3_1 _16562_ (.A(_09059_),
    .B(_08470_),
    .C(_08546_),
    .X(_09205_));
 sky130_fd_sc_hd__a21boi_1 _16563_ (.A1(_09089_),
    .A2(_09205_),
    .B1_N(_09192_),
    .Y(_09206_));
 sky130_fd_sc_hd__a31o_4 _16564_ (.A1(_08549_),
    .A2(_08957_),
    .A3(_09204_),
    .B1(_09206_),
    .X(_09207_));
 sky130_fd_sc_hd__nor2_1 _16565_ (.A(_09188_),
    .B(_09191_),
    .Y(_09208_));
 sky130_fd_sc_hd__o21ai_1 _16566_ (.A1(_09175_),
    .A2(_09176_),
    .B1(_09178_),
    .Y(_09209_));
 sky130_fd_sc_hd__a21o_1 _16567_ (.A1(_09090_),
    .A2(_09112_),
    .B1(_09110_),
    .X(_09210_));
 sky130_fd_sc_hd__nor2_1 _16568_ (.A(_08054_),
    .B(_09029_),
    .Y(_09211_));
 sky130_fd_sc_hd__or3b_1 _16569_ (.A(_08160_),
    .B(_09165_),
    .C_N(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__a31o_1 _16570_ (.A1(\rbzero.wall_tracer.visualWallDist[7] ),
    .A2(_04015_),
    .A3(_08416_),
    .B1(_09211_),
    .X(_09213_));
 sky130_fd_sc_hd__nand2_1 _16571_ (.A(_09212_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__nand2_4 _16572_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_04015_),
    .Y(_09215_));
 sky130_fd_sc_hd__or2_1 _16573_ (.A(_05210_),
    .B(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__clkbuf_4 _16574_ (.A(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__nor2_1 _16575_ (.A(_08162_),
    .B(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__xnor2_1 _16576_ (.A(_09214_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(_09161_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__or2_1 _16578_ (.A(_09161_),
    .B(_09219_),
    .X(_09221_));
 sky130_fd_sc_hd__and2_1 _16579_ (.A(_09220_),
    .B(_09221_),
    .X(_09222_));
 sky130_fd_sc_hd__a21bo_1 _16580_ (.A1(_09170_),
    .A2(_09172_),
    .B1_N(_09169_),
    .X(_09223_));
 sky130_fd_sc_hd__nand2_1 _16581_ (.A(_09092_),
    .B(_09095_),
    .Y(_09224_));
 sky130_fd_sc_hd__or3_1 _16582_ (.A(_08821_),
    .B(_08823_),
    .C(_08419_),
    .X(_09225_));
 sky130_fd_sc_hd__o22ai_1 _16583_ (.A1(_08823_),
    .A2(_08159_),
    .B1(_08151_),
    .B2(_09096_),
    .Y(_09226_));
 sky130_fd_sc_hd__nand2_1 _16584_ (.A(_09225_),
    .B(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__nor2_1 _16585_ (.A(_08329_),
    .B(_08427_),
    .Y(_09228_));
 sky130_fd_sc_hd__xor2_1 _16586_ (.A(_09227_),
    .B(_09228_),
    .X(_09229_));
 sky130_fd_sc_hd__xnor2_1 _16587_ (.A(_09224_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__xnor2_1 _16588_ (.A(_09223_),
    .B(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__a21oi_1 _16589_ (.A1(_09003_),
    .A2(_09006_),
    .B1(_09173_),
    .Y(_09232_));
 sky130_fd_sc_hd__a21oi_1 _16590_ (.A1(_09167_),
    .A2(_09174_),
    .B1(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__nor2_1 _16591_ (.A(_09231_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__and2_1 _16592_ (.A(_09231_),
    .B(_09233_),
    .X(_09235_));
 sky130_fd_sc_hd__nor2_1 _16593_ (.A(_09234_),
    .B(_09235_),
    .Y(_09236_));
 sky130_fd_sc_hd__xor2_1 _16594_ (.A(_09222_),
    .B(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__xnor2_1 _16595_ (.A(_09210_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__xnor2_1 _16596_ (.A(_09209_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__a21o_1 _16597_ (.A1(_09098_),
    .A2(_09108_),
    .B1(_09106_),
    .X(_09240_));
 sky130_fd_sc_hd__nand2_1 _16598_ (.A(_09118_),
    .B(_09123_),
    .Y(_09241_));
 sky130_fd_sc_hd__or2b_1 _16599_ (.A(_09124_),
    .B_N(_09116_),
    .X(_09242_));
 sky130_fd_sc_hd__buf_2 _16600_ (.A(_08075_),
    .X(_09243_));
 sky130_fd_sc_hd__or4_1 _16601_ (.A(_07932_),
    .B(_07938_),
    .C(_08035_),
    .D(_08046_),
    .X(_09244_));
 sky130_fd_sc_hd__buf_2 _16602_ (.A(_07938_),
    .X(_09245_));
 sky130_fd_sc_hd__o22ai_1 _16603_ (.A1(_07932_),
    .A2(_08129_),
    .B1(_08047_),
    .B2(_09245_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(_09244_),
    .B(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__or3_1 _16605_ (.A(_09243_),
    .B(_08059_),
    .C(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__clkbuf_4 _16606_ (.A(_09243_),
    .X(_09249_));
 sky130_fd_sc_hd__o21ai_1 _16607_ (.A1(_09249_),
    .A2(_08356_),
    .B1(_09247_),
    .Y(_09250_));
 sky130_fd_sc_hd__and2_1 _16608_ (.A(_09248_),
    .B(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__or4_1 _16609_ (.A(_08282_),
    .B(_08383_),
    .C(_08111_),
    .D(_08570_),
    .X(_09252_));
 sky130_fd_sc_hd__o22ai_1 _16610_ (.A1(_08383_),
    .A2(_08111_),
    .B1(_08570_),
    .B2(_08282_),
    .Y(_09253_));
 sky130_fd_sc_hd__nand2_1 _16611_ (.A(_09252_),
    .B(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__or2_1 _16612_ (.A(_07996_),
    .B(_09103_),
    .X(_09255_));
 sky130_fd_sc_hd__xnor2_1 _16613_ (.A(_09254_),
    .B(_09255_),
    .Y(_09256_));
 sky130_fd_sc_hd__nand2_1 _16614_ (.A(_09009_),
    .B(_09099_),
    .Y(_09257_));
 sky130_fd_sc_hd__o31a_1 _16615_ (.A1(_07932_),
    .A2(_09103_),
    .A3(_09100_),
    .B1(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__nor2_1 _16616_ (.A(_09256_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__and2_1 _16617_ (.A(_09256_),
    .B(_09258_),
    .X(_09260_));
 sky130_fd_sc_hd__nor2_1 _16618_ (.A(_09259_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__xnor2_1 _16619_ (.A(_09251_),
    .B(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__a21o_1 _16620_ (.A1(_09241_),
    .A2(_09242_),
    .B1(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__nand3_1 _16621_ (.A(_09241_),
    .B(_09242_),
    .C(_09262_),
    .Y(_09264_));
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(_09263_),
    .B(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__xnor2_1 _16623_ (.A(_09240_),
    .B(_09265_),
    .Y(_09266_));
 sky130_fd_sc_hd__or3_1 _16624_ (.A(_08383_),
    .B(_09114_),
    .C(_09121_),
    .X(_09267_));
 sky130_fd_sc_hd__a21bo_1 _16625_ (.A1(_08963_),
    .A2(_09119_),
    .B1_N(_09267_),
    .X(_09268_));
 sky130_fd_sc_hd__a22o_1 _16626_ (.A1(_09128_),
    .A2(_09130_),
    .B1(_09131_),
    .B2(_09127_),
    .X(_09269_));
 sky130_fd_sc_hd__nor2_1 _16627_ (.A(_08283_),
    .B(_08189_),
    .Y(_09270_));
 sky130_fd_sc_hd__xnor2_1 _16628_ (.A(_09119_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__nor2_1 _16629_ (.A(_09114_),
    .B(_08204_),
    .Y(_09272_));
 sky130_fd_sc_hd__xnor2_1 _16630_ (.A(_09271_),
    .B(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__xnor2_1 _16631_ (.A(_09269_),
    .B(_09273_),
    .Y(_09274_));
 sky130_fd_sc_hd__xnor2_1 _16632_ (.A(_09268_),
    .B(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__clkbuf_4 _16633_ (.A(_08971_),
    .X(_09276_));
 sky130_fd_sc_hd__nor2_1 _16634_ (.A(_09117_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__a21oi_1 _16635_ (.A1(_08242_),
    .A2(_09129_),
    .B1(_08180_),
    .Y(_09278_));
 sky130_fd_sc_hd__nand2_2 _16636_ (.A(_05209_),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_09279_));
 sky130_fd_sc_hd__a21oi_1 _16637_ (.A1(_08237_),
    .A2(_09279_),
    .B1(_08170_),
    .Y(_09280_));
 sky130_fd_sc_hd__xor2_1 _16638_ (.A(_09278_),
    .B(_09280_),
    .X(_09281_));
 sky130_fd_sc_hd__xor2_1 _16639_ (.A(_09277_),
    .B(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__buf_6 _16640_ (.A(_08230_),
    .X(_09283_));
 sky130_fd_sc_hd__nand2_1 _16641_ (.A(_09283_),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_09284_));
 sky130_fd_sc_hd__o21ai_1 _16642_ (.A1(_07575_),
    .A2(_08983_),
    .B1(_07579_),
    .Y(_09285_));
 sky130_fd_sc_hd__or3_1 _16643_ (.A(_07575_),
    .B(_07579_),
    .C(_08983_),
    .X(_09286_));
 sky130_fd_sc_hd__a31o_1 _16644_ (.A1(_05194_),
    .A2(_09285_),
    .A3(_09286_),
    .B1(_08224_),
    .X(_09287_));
 sky130_fd_sc_hd__a21o_1 _16645_ (.A1(_09284_),
    .A2(_09287_),
    .B1(_05210_),
    .X(_09288_));
 sky130_fd_sc_hd__o22ai_1 _16646_ (.A1(_08215_),
    .A2(_08985_),
    .B1(_09138_),
    .B2(_08519_),
    .Y(_09289_));
 sky130_fd_sc_hd__or4_1 _16647_ (.A(_08215_),
    .B(_08519_),
    .C(_08985_),
    .D(_09138_),
    .X(_09290_));
 sky130_fd_sc_hd__or4bb_1 _16648_ (.A(_08239_),
    .B(_09288_),
    .C_N(_09289_),
    .D_N(_09290_),
    .X(_09291_));
 sky130_fd_sc_hd__buf_4 _16649_ (.A(_09288_),
    .X(_09292_));
 sky130_fd_sc_hd__a2bb2o_1 _16650_ (.A1_N(_08239_),
    .A2_N(_09292_),
    .B1(_09289_),
    .B2(_09290_),
    .X(_09293_));
 sky130_fd_sc_hd__or2_2 _16651_ (.A(_05211_),
    .B(_09138_),
    .X(_09294_));
 sky130_fd_sc_hd__or2_1 _16652_ (.A(_09133_),
    .B(_09134_),
    .X(_09295_));
 sky130_fd_sc_hd__o31ai_1 _16653_ (.A1(_08239_),
    .A2(_09135_),
    .A3(_09294_),
    .B1(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__nand3_1 _16654_ (.A(_09291_),
    .B(_09293_),
    .C(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__a21o_1 _16655_ (.A1(_09291_),
    .A2(_09293_),
    .B1(_09296_),
    .X(_09298_));
 sky130_fd_sc_hd__nand3_1 _16656_ (.A(_09282_),
    .B(_09297_),
    .C(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__a21o_1 _16657_ (.A1(_09297_),
    .A2(_09298_),
    .B1(_09282_),
    .X(_09300_));
 sky130_fd_sc_hd__or2b_1 _16658_ (.A(_09143_),
    .B_N(_09140_),
    .X(_09301_));
 sky130_fd_sc_hd__a21bo_1 _16659_ (.A1(_09132_),
    .A2(_09144_),
    .B1_N(_09301_),
    .X(_09302_));
 sky130_fd_sc_hd__nand3_1 _16660_ (.A(_09299_),
    .B(_09300_),
    .C(_09302_),
    .Y(_09303_));
 sky130_fd_sc_hd__a21o_1 _16661_ (.A1(_09299_),
    .A2(_09300_),
    .B1(_09302_),
    .X(_09304_));
 sky130_fd_sc_hd__nand3_1 _16662_ (.A(_09275_),
    .B(_09303_),
    .C(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__a21o_1 _16663_ (.A1(_09303_),
    .A2(_09304_),
    .B1(_09275_),
    .X(_09306_));
 sky130_fd_sc_hd__nor2_1 _16664_ (.A(_09145_),
    .B(_09147_),
    .Y(_09307_));
 sky130_fd_sc_hd__a21o_1 _16665_ (.A1(_09125_),
    .A2(_09148_),
    .B1(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__nand3_1 _16666_ (.A(_09305_),
    .B(_09306_),
    .C(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__a21o_1 _16667_ (.A1(_09305_),
    .A2(_09306_),
    .B1(_09308_),
    .X(_09310_));
 sky130_fd_sc_hd__nand3_1 _16668_ (.A(_09266_),
    .B(_09309_),
    .C(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__a21o_1 _16669_ (.A1(_09309_),
    .A2(_09310_),
    .B1(_09266_),
    .X(_09312_));
 sky130_fd_sc_hd__and2b_1 _16670_ (.A_N(_09149_),
    .B(_09151_),
    .X(_09313_));
 sky130_fd_sc_hd__a21o_1 _16671_ (.A1(_09113_),
    .A2(_09152_),
    .B1(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__and3_1 _16672_ (.A(_09311_),
    .B(_09312_),
    .C(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__a21oi_1 _16673_ (.A1(_09311_),
    .A2(_09312_),
    .B1(_09314_),
    .Y(_09316_));
 sky130_fd_sc_hd__nor2_1 _16674_ (.A(_09315_),
    .B(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__xnor2_1 _16675_ (.A(_09239_),
    .B(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__nor2_1 _16676_ (.A(_09153_),
    .B(_09155_),
    .Y(_09319_));
 sky130_fd_sc_hd__a21oi_1 _16677_ (.A1(_09156_),
    .A2(_09182_),
    .B1(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__xnor2_1 _16678_ (.A(_09318_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__or2b_1 _16679_ (.A(_09181_),
    .B_N(_09158_),
    .X(_09322_));
 sky130_fd_sc_hd__a21boi_1 _16680_ (.A1(_09160_),
    .A2(_09180_),
    .B1_N(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__xnor2_1 _16681_ (.A(_09321_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__or2_1 _16682_ (.A(_09183_),
    .B(_09185_),
    .X(_09325_));
 sky130_fd_sc_hd__o21a_1 _16683_ (.A1(_09186_),
    .A2(_09187_),
    .B1(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__xor2_1 _16684_ (.A(_09324_),
    .B(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__nand2_1 _16685_ (.A(_09208_),
    .B(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__or2_1 _16686_ (.A(_09208_),
    .B(_09327_),
    .X(_09329_));
 sky130_fd_sc_hd__and2_2 _16687_ (.A(_09328_),
    .B(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__xnor2_4 _16688_ (.A(_09207_),
    .B(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__inv_2 _16689_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_09332_));
 sky130_fd_sc_hd__mux2_1 _16690_ (.A0(_09332_),
    .A1(_07949_),
    .S(_07895_),
    .X(_09333_));
 sky130_fd_sc_hd__nor2_1 _16691_ (.A(_09331_),
    .B(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _16692_ (.A(_09331_),
    .B(_09333_),
    .Y(_09335_));
 sky130_fd_sc_hd__or2b_1 _16693_ (.A(_09334_),
    .B_N(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__a21o_1 _16694_ (.A1(_09198_),
    .A2(_09200_),
    .B1(_09197_),
    .X(_09337_));
 sky130_fd_sc_hd__xnor2_1 _16695_ (.A(_09336_),
    .B(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__xnor2_1 _16696_ (.A(_09082_),
    .B(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__or2_1 _16697_ (.A(\rbzero.wall_tracer.texu[2] ),
    .B(_09085_),
    .X(_09340_));
 sky130_fd_sc_hd__o211a_1 _16698_ (.A1(_05194_),
    .A2(_09339_),
    .B1(_09340_),
    .C1(_07642_),
    .X(_00513_));
 sky130_fd_sc_hd__a21bo_1 _16699_ (.A1(_09207_),
    .A2(_09330_),
    .B1_N(_09328_),
    .X(_09341_));
 sky130_fd_sc_hd__or2_2 _16700_ (.A(_09324_),
    .B(_09326_),
    .X(_09342_));
 sky130_fd_sc_hd__or2b_1 _16701_ (.A(_09238_),
    .B_N(_09209_),
    .X(_09343_));
 sky130_fd_sc_hd__a21boi_1 _16702_ (.A1(_09210_),
    .A2(_09237_),
    .B1_N(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__nor2_1 _16703_ (.A(_09220_),
    .B(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__and2_1 _16704_ (.A(_09220_),
    .B(_09344_),
    .X(_09346_));
 sky130_fd_sc_hd__nor2_1 _16705_ (.A(_09345_),
    .B(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__a21o_1 _16706_ (.A1(_09222_),
    .A2(_09236_),
    .B1(_09234_),
    .X(_09348_));
 sky130_fd_sc_hd__or2b_1 _16707_ (.A(_09265_),
    .B_N(_09240_),
    .X(_09349_));
 sky130_fd_sc_hd__nand2_4 _16708_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_04015_),
    .Y(_09350_));
 sky130_fd_sc_hd__or2_1 _16709_ (.A(_05210_),
    .B(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__or2_1 _16710_ (.A(_08162_),
    .B(_09351_),
    .X(_09352_));
 sky130_fd_sc_hd__inv_2 _16711_ (.A(_09028_),
    .Y(_09353_));
 sky130_fd_sc_hd__nand2_1 _16712_ (.A(_08331_),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__nor2_1 _16713_ (.A(_08054_),
    .B(_09164_),
    .Y(_09355_));
 sky130_fd_sc_hd__xnor2_1 _16714_ (.A(_09354_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__nor2_1 _16715_ (.A(_08062_),
    .B(_09217_),
    .Y(_09357_));
 sky130_fd_sc_hd__xnor2_1 _16716_ (.A(_09356_),
    .B(_09357_),
    .Y(_09358_));
 sky130_fd_sc_hd__clkbuf_4 _16717_ (.A(_09217_),
    .X(_09359_));
 sky130_fd_sc_hd__o31a_1 _16718_ (.A1(_08162_),
    .A2(_09214_),
    .A3(_09359_),
    .B1(_09212_),
    .X(_09360_));
 sky130_fd_sc_hd__xor2_1 _16719_ (.A(_09358_),
    .B(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__xnor2_1 _16720_ (.A(_09352_),
    .B(_09361_),
    .Y(_09362_));
 sky130_fd_sc_hd__a21bo_1 _16721_ (.A1(_09226_),
    .A2(_09228_),
    .B1_N(_09225_),
    .X(_09363_));
 sky130_fd_sc_hd__nand2_1 _16722_ (.A(_09244_),
    .B(_09248_),
    .Y(_09364_));
 sky130_fd_sc_hd__or3_1 _16723_ (.A(_09243_),
    .B(_08821_),
    .C(_08419_),
    .X(_09365_));
 sky130_fd_sc_hd__o22ai_1 _16724_ (.A1(_08821_),
    .A2(_08159_),
    .B1(_08151_),
    .B2(_09243_),
    .Y(_09366_));
 sky130_fd_sc_hd__nand2_1 _16725_ (.A(_09365_),
    .B(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__buf_2 _16726_ (.A(_08823_),
    .X(_09368_));
 sky130_fd_sc_hd__nor2_1 _16727_ (.A(_09368_),
    .B(_08427_),
    .Y(_09369_));
 sky130_fd_sc_hd__xor2_1 _16728_ (.A(_09367_),
    .B(_09369_),
    .X(_09370_));
 sky130_fd_sc_hd__xnor2_1 _16729_ (.A(_09364_),
    .B(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__xnor2_1 _16730_ (.A(_09363_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__a21oi_1 _16731_ (.A1(_09092_),
    .A2(_09095_),
    .B1(_09229_),
    .Y(_09373_));
 sky130_fd_sc_hd__a21oi_1 _16732_ (.A1(_09223_),
    .A2(_09230_),
    .B1(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_1 _16733_ (.A(_09372_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__and2_1 _16734_ (.A(_09372_),
    .B(_09374_),
    .X(_09376_));
 sky130_fd_sc_hd__nor2_1 _16735_ (.A(_09375_),
    .B(_09376_),
    .Y(_09377_));
 sky130_fd_sc_hd__xnor2_1 _16736_ (.A(_09362_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__a21o_1 _16737_ (.A1(_09263_),
    .A2(_09349_),
    .B1(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__nand3_1 _16738_ (.A(_09263_),
    .B(_09349_),
    .C(_09378_),
    .Y(_09380_));
 sky130_fd_sc_hd__nand2_1 _16739_ (.A(_09379_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__xnor2_1 _16740_ (.A(_09348_),
    .B(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__a21o_1 _16741_ (.A1(_09251_),
    .A2(_09261_),
    .B1(_09259_),
    .X(_09383_));
 sky130_fd_sc_hd__or2_1 _16742_ (.A(_09269_),
    .B(_09273_),
    .X(_09384_));
 sky130_fd_sc_hd__and2_1 _16743_ (.A(_09269_),
    .B(_09273_),
    .X(_09385_));
 sky130_fd_sc_hd__a21o_1 _16744_ (.A1(_09268_),
    .A2(_09384_),
    .B1(_09385_),
    .X(_09386_));
 sky130_fd_sc_hd__or4_1 _16745_ (.A(_07996_),
    .B(_08705_),
    .C(_08035_),
    .D(_08046_),
    .X(_09387_));
 sky130_fd_sc_hd__o22ai_1 _16746_ (.A1(_07996_),
    .A2(_08129_),
    .B1(_08047_),
    .B2(_08705_),
    .Y(_09388_));
 sky130_fd_sc_hd__nand2_1 _16747_ (.A(_09387_),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__or3_1 _16748_ (.A(_09245_),
    .B(_08059_),
    .C(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__clkbuf_4 _16749_ (.A(_09245_),
    .X(_09391_));
 sky130_fd_sc_hd__o21ai_1 _16750_ (.A1(_09391_),
    .A2(_08356_),
    .B1(_09389_),
    .Y(_09392_));
 sky130_fd_sc_hd__and2_1 _16751_ (.A(_09390_),
    .B(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__or2_1 _16752_ (.A(_09254_),
    .B(_09255_),
    .X(_09394_));
 sky130_fd_sc_hd__nor2_1 _16753_ (.A(_08383_),
    .B(_08570_),
    .Y(_09395_));
 sky130_fd_sc_hd__and2b_1 _16754_ (.A_N(_08111_),
    .B(_08264_),
    .X(_09396_));
 sky130_fd_sc_hd__xnor2_1 _16755_ (.A(_09395_),
    .B(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__or2_1 _16756_ (.A(_08282_),
    .B(_09103_),
    .X(_09398_));
 sky130_fd_sc_hd__xnor2_1 _16757_ (.A(_09397_),
    .B(_09398_),
    .Y(_09399_));
 sky130_fd_sc_hd__a21oi_1 _16758_ (.A1(_09252_),
    .A2(_09394_),
    .B1(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__and3_1 _16759_ (.A(_09252_),
    .B(_09394_),
    .C(_09399_),
    .X(_09401_));
 sky130_fd_sc_hd__nor2_1 _16760_ (.A(_09400_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__xnor2_1 _16761_ (.A(_09393_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__xor2_1 _16762_ (.A(_09386_),
    .B(_09403_),
    .X(_09404_));
 sky130_fd_sc_hd__xnor2_1 _16763_ (.A(_09383_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__or3_1 _16764_ (.A(_09114_),
    .B(_08204_),
    .C(_09271_),
    .X(_09406_));
 sky130_fd_sc_hd__a21bo_1 _16765_ (.A1(_09119_),
    .A2(_09270_),
    .B1_N(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__a22oi_2 _16766_ (.A1(_09278_),
    .A2(_09280_),
    .B1(_09281_),
    .B2(_09277_),
    .Y(_09408_));
 sky130_fd_sc_hd__nor2_1 _16767_ (.A(_08284_),
    .B(_09276_),
    .Y(_09409_));
 sky130_fd_sc_hd__o22a_1 _16768_ (.A1(_08284_),
    .A2(_09126_),
    .B1(_09276_),
    .B2(_08283_),
    .X(_09410_));
 sky130_fd_sc_hd__a21o_1 _16769_ (.A1(_09270_),
    .A2(_09409_),
    .B1(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__or2_1 _16770_ (.A(_09114_),
    .B(_08178_),
    .X(_09412_));
 sky130_fd_sc_hd__xor2_2 _16771_ (.A(_09411_),
    .B(_09412_),
    .X(_09413_));
 sky130_fd_sc_hd__xnor2_2 _16772_ (.A(_09408_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__xor2_2 _16773_ (.A(_09407_),
    .B(_09414_),
    .X(_09415_));
 sky130_fd_sc_hd__and2_1 _16774_ (.A(_08242_),
    .B(_09129_),
    .X(_09416_));
 sky130_fd_sc_hd__clkbuf_4 _16775_ (.A(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__nor2_1 _16776_ (.A(_09117_),
    .B(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__a21o_1 _16777_ (.A1(_08237_),
    .A2(_09279_),
    .B1(_08180_),
    .X(_09419_));
 sky130_fd_sc_hd__nand2_1 _16778_ (.A(_05210_),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_09420_));
 sky130_fd_sc_hd__a21oi_1 _16779_ (.A1(_09141_),
    .A2(_09420_),
    .B1(_08170_),
    .Y(_09421_));
 sky130_fd_sc_hd__xnor2_1 _16780_ (.A(_09419_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__and2_1 _16781_ (.A(_09418_),
    .B(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__nor2_1 _16782_ (.A(_09418_),
    .B(_09422_),
    .Y(_09424_));
 sky130_fd_sc_hd__nor2_1 _16783_ (.A(_09423_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__nor2_1 _16784_ (.A(_08377_),
    .B(_09138_),
    .Y(_09426_));
 sky130_fd_sc_hd__or4_1 _16785_ (.A(_07598_),
    .B(_09283_),
    .C(_05209_),
    .D(_09287_),
    .X(_09427_));
 sky130_fd_sc_hd__xnor2_2 _16786_ (.A(_09426_),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand2_1 _16787_ (.A(_08230_),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_09429_));
 sky130_fd_sc_hd__or2_1 _16788_ (.A(_07579_),
    .B(_07582_),
    .X(_09430_));
 sky130_fd_sc_hd__nor3_2 _16789_ (.A(_07575_),
    .B(_08983_),
    .C(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__o31a_1 _16790_ (.A1(_07575_),
    .A2(_07579_),
    .A3(_08983_),
    .B1(_07582_),
    .X(_09432_));
 sky130_fd_sc_hd__o31ai_4 _16791_ (.A1(_09085_),
    .A2(_09431_),
    .A3(_09432_),
    .B1(_08235_),
    .Y(_09433_));
 sky130_fd_sc_hd__a21o_2 _16792_ (.A1(_09429_),
    .A2(_09433_),
    .B1(_05209_),
    .X(_09434_));
 sky130_fd_sc_hd__nor2_1 _16793_ (.A(_08239_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__xnor2_2 _16794_ (.A(_09428_),
    .B(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__nand2_1 _16795_ (.A(_09290_),
    .B(_09291_),
    .Y(_09437_));
 sky130_fd_sc_hd__xnor2_2 _16796_ (.A(_09436_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__xnor2_2 _16797_ (.A(_09425_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__and2_1 _16798_ (.A(_09297_),
    .B(_09299_),
    .X(_09440_));
 sky130_fd_sc_hd__xor2_2 _16799_ (.A(_09439_),
    .B(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__xnor2_2 _16800_ (.A(_09415_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__and2_1 _16801_ (.A(_09303_),
    .B(_09305_),
    .X(_09443_));
 sky130_fd_sc_hd__xor2_1 _16802_ (.A(_09442_),
    .B(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__xnor2_1 _16803_ (.A(_09405_),
    .B(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__and2_1 _16804_ (.A(_09309_),
    .B(_09311_),
    .X(_09446_));
 sky130_fd_sc_hd__xor2_1 _16805_ (.A(_09445_),
    .B(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__xnor2_1 _16806_ (.A(_09382_),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__a21oi_1 _16807_ (.A1(_09239_),
    .A2(_09317_),
    .B1(_09315_),
    .Y(_09449_));
 sky130_fd_sc_hd__xor2_1 _16808_ (.A(_09448_),
    .B(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__xnor2_1 _16809_ (.A(_09347_),
    .B(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__or2_1 _16810_ (.A(_09318_),
    .B(_09320_),
    .X(_09452_));
 sky130_fd_sc_hd__o21a_1 _16811_ (.A1(_09321_),
    .A2(_09323_),
    .B1(_09452_),
    .X(_09453_));
 sky130_fd_sc_hd__nor2_1 _16812_ (.A(_09451_),
    .B(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__and2_1 _16813_ (.A(_09451_),
    .B(_09453_),
    .X(_09455_));
 sky130_fd_sc_hd__or2_2 _16814_ (.A(_09454_),
    .B(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__xor2_4 _16815_ (.A(_09342_),
    .B(_09456_),
    .X(_09457_));
 sky130_fd_sc_hd__xnor2_4 _16816_ (.A(_09341_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__clkinv_2 _16817_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_09459_));
 sky130_fd_sc_hd__mux2_1 _16818_ (.A0(_09459_),
    .A1(_08067_),
    .S(_07895_),
    .X(_09460_));
 sky130_fd_sc_hd__nor2_1 _16819_ (.A(_09458_),
    .B(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__and2_1 _16820_ (.A(_09458_),
    .B(_09460_),
    .X(_09462_));
 sky130_fd_sc_hd__or2_1 _16821_ (.A(_09461_),
    .B(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__a21oi_1 _16822_ (.A1(_09335_),
    .A2(_09337_),
    .B1(_09334_),
    .Y(_09464_));
 sky130_fd_sc_hd__nor2_1 _16823_ (.A(_09463_),
    .B(_09464_),
    .Y(_09465_));
 sky130_fd_sc_hd__and2_1 _16824_ (.A(_09463_),
    .B(_09464_),
    .X(_09466_));
 sky130_fd_sc_hd__nor2_1 _16825_ (.A(_09465_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__nor2_1 _16826_ (.A(_09082_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__a21o_1 _16827_ (.A1(_09082_),
    .A2(_09467_),
    .B1(_05194_),
    .X(_09469_));
 sky130_fd_sc_hd__o221a_1 _16828_ (.A1(\rbzero.wall_tracer.texu[3] ),
    .A2(_09085_),
    .B1(_09468_),
    .B2(_09469_),
    .C1(_07642_),
    .X(_00514_));
 sky130_fd_sc_hd__or2_1 _16829_ (.A(_09461_),
    .B(_09465_),
    .X(_09470_));
 sky130_fd_sc_hd__or2b_1 _16830_ (.A(_09381_),
    .B_N(_09348_),
    .X(_09471_));
 sky130_fd_sc_hd__or2b_1 _16831_ (.A(_09352_),
    .B_N(_09361_),
    .X(_09472_));
 sky130_fd_sc_hd__o21a_1 _16832_ (.A1(_09358_),
    .A2(_09360_),
    .B1(_09472_),
    .X(_09473_));
 sky130_fd_sc_hd__a21oi_2 _16833_ (.A1(_09379_),
    .A2(_09471_),
    .B1(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__and3_1 _16834_ (.A(_09379_),
    .B(_09471_),
    .C(_09473_),
    .X(_09475_));
 sky130_fd_sc_hd__nor2_1 _16835_ (.A(_09474_),
    .B(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__a21o_1 _16836_ (.A1(_09362_),
    .A2(_09377_),
    .B1(_09375_),
    .X(_09477_));
 sky130_fd_sc_hd__or2b_1 _16837_ (.A(_09403_),
    .B_N(_09386_),
    .X(_09478_));
 sky130_fd_sc_hd__or2b_1 _16838_ (.A(_09404_),
    .B_N(_09383_),
    .X(_09479_));
 sky130_fd_sc_hd__clkbuf_4 _16839_ (.A(_09351_),
    .X(_09480_));
 sky130_fd_sc_hd__nand2_2 _16840_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_04015_),
    .Y(_09481_));
 sky130_fd_sc_hd__or2_1 _16841_ (.A(_05211_),
    .B(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__buf_2 _16842_ (.A(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__clkbuf_4 _16843_ (.A(_09483_),
    .X(_09484_));
 sky130_fd_sc_hd__o22ai_1 _16844_ (.A1(_08160_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_08162_),
    .Y(_09485_));
 sky130_fd_sc_hd__or3_1 _16845_ (.A(_08160_),
    .B(_09352_),
    .C(_09484_),
    .X(_09486_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(_09485_),
    .B(_09486_),
    .Y(_09487_));
 sky130_fd_sc_hd__nor2_1 _16847_ (.A(_08054_),
    .B(_09216_),
    .Y(_09488_));
 sky130_fd_sc_hd__o22a_1 _16848_ (.A1(_08823_),
    .A2(_09028_),
    .B1(_09164_),
    .B2(_08329_),
    .X(_09489_));
 sky130_fd_sc_hd__or3_1 _16849_ (.A(_08823_),
    .B(_09164_),
    .C(_09354_),
    .X(_09490_));
 sky130_fd_sc_hd__and2b_1 _16850_ (.A_N(_09489_),
    .B(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__xnor2_1 _16851_ (.A(_09488_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(_09356_),
    .B(_09357_),
    .Y(_09493_));
 sky130_fd_sc_hd__o31a_1 _16853_ (.A1(_08335_),
    .A2(_09165_),
    .A3(_09354_),
    .B1(_09493_),
    .X(_09494_));
 sky130_fd_sc_hd__nor2_1 _16854_ (.A(_09492_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__and2_1 _16855_ (.A(_09492_),
    .B(_09494_),
    .X(_09496_));
 sky130_fd_sc_hd__nor2_1 _16856_ (.A(_09495_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__xnor2_1 _16857_ (.A(_09487_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__a21bo_1 _16858_ (.A1(_09366_),
    .A2(_09369_),
    .B1_N(_09365_),
    .X(_09499_));
 sky130_fd_sc_hd__nand2_1 _16859_ (.A(_09387_),
    .B(_09390_),
    .Y(_09500_));
 sky130_fd_sc_hd__nor2_1 _16860_ (.A(_09096_),
    .B(_08427_),
    .Y(_09501_));
 sky130_fd_sc_hd__o22a_1 _16861_ (.A1(_09243_),
    .A2(_08159_),
    .B1(_08150_),
    .B2(_09245_),
    .X(_09502_));
 sky130_fd_sc_hd__or4_1 _16862_ (.A(_09245_),
    .B(_08075_),
    .C(_08159_),
    .D(_08150_),
    .X(_09503_));
 sky130_fd_sc_hd__and2b_1 _16863_ (.A_N(_09502_),
    .B(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__xnor2_1 _16864_ (.A(_09501_),
    .B(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__xnor2_1 _16865_ (.A(_09500_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__xnor2_1 _16866_ (.A(_09499_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__a21oi_1 _16867_ (.A1(_09244_),
    .A2(_09248_),
    .B1(_09370_),
    .Y(_09508_));
 sky130_fd_sc_hd__a21oi_1 _16868_ (.A1(_09363_),
    .A2(_09371_),
    .B1(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__nor2_1 _16869_ (.A(_09507_),
    .B(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__and2_1 _16870_ (.A(_09507_),
    .B(_09509_),
    .X(_09511_));
 sky130_fd_sc_hd__nor2_1 _16871_ (.A(_09510_),
    .B(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__xnor2_1 _16872_ (.A(_09498_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__a21o_1 _16873_ (.A1(_09478_),
    .A2(_09479_),
    .B1(_09513_),
    .X(_09514_));
 sky130_fd_sc_hd__nand3_1 _16874_ (.A(_09478_),
    .B(_09479_),
    .C(_09513_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_1 _16875_ (.A(_09514_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__xnor2_1 _16876_ (.A(_09477_),
    .B(_09516_),
    .Y(_09517_));
 sky130_fd_sc_hd__a21o_1 _16877_ (.A1(_09393_),
    .A2(_09402_),
    .B1(_09400_),
    .X(_09518_));
 sky130_fd_sc_hd__and2b_1 _16878_ (.A_N(_09408_),
    .B(_09413_),
    .X(_09519_));
 sky130_fd_sc_hd__a21o_1 _16879_ (.A1(_09407_),
    .A2(_09414_),
    .B1(_09519_),
    .X(_09520_));
 sky130_fd_sc_hd__or4_1 _16880_ (.A(_08282_),
    .B(_07994_),
    .C(_08035_),
    .D(_08046_),
    .X(_09521_));
 sky130_fd_sc_hd__buf_2 _16881_ (.A(_07994_),
    .X(_09522_));
 sky130_fd_sc_hd__o22ai_1 _16882_ (.A1(_08282_),
    .A2(_08129_),
    .B1(_08047_),
    .B2(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__nand2_1 _16883_ (.A(_09521_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__or3_1 _16884_ (.A(_08705_),
    .B(_08059_),
    .C(_09524_),
    .X(_09525_));
 sky130_fd_sc_hd__clkbuf_4 _16885_ (.A(_08705_),
    .X(_09526_));
 sky130_fd_sc_hd__o21ai_1 _16886_ (.A1(_09526_),
    .A2(_08356_),
    .B1(_09524_),
    .Y(_09527_));
 sky130_fd_sc_hd__and2_1 _16887_ (.A(_09525_),
    .B(_09527_),
    .X(_09528_));
 sky130_fd_sc_hd__nor2_1 _16888_ (.A(_08204_),
    .B(_08570_),
    .Y(_09529_));
 sky130_fd_sc_hd__nor2_1 _16889_ (.A(_08178_),
    .B(_08111_),
    .Y(_09530_));
 sky130_fd_sc_hd__xnor2_2 _16890_ (.A(_09529_),
    .B(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__or2_1 _16891_ (.A(_08383_),
    .B(_09103_),
    .X(_09532_));
 sky130_fd_sc_hd__xnor2_2 _16892_ (.A(_09531_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__o2bb2a_1 _16893_ (.A1_N(_09395_),
    .A2_N(_09396_),
    .B1(_09397_),
    .B2(_09398_),
    .X(_09534_));
 sky130_fd_sc_hd__xor2_2 _16894_ (.A(_09533_),
    .B(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__xnor2_2 _16895_ (.A(_09528_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__xor2_1 _16896_ (.A(_09520_),
    .B(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__xnor2_1 _16897_ (.A(_09518_),
    .B(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__a2bb2o_1 _16898_ (.A1_N(_09410_),
    .A2_N(_09412_),
    .B1(_09270_),
    .B2(_09409_),
    .X(_09539_));
 sky130_fd_sc_hd__and2_1 _16899_ (.A(_08985_),
    .B(_09420_),
    .X(_09540_));
 sky130_fd_sc_hd__or3_1 _16900_ (.A(_08170_),
    .B(_09419_),
    .C(_09540_),
    .X(_09541_));
 sky130_fd_sc_hd__inv_2 _16901_ (.A(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__a21oi_1 _16902_ (.A1(_08242_),
    .A2(_09129_),
    .B1(_08283_),
    .Y(_09543_));
 sky130_fd_sc_hd__xnor2_1 _16903_ (.A(_09409_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nor2_2 _16904_ (.A(_07959_),
    .B(_09126_),
    .Y(_09545_));
 sky130_fd_sc_hd__xnor2_1 _16905_ (.A(_09544_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__o21a_1 _16906_ (.A1(_09542_),
    .A2(_09423_),
    .B1(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__a211o_1 _16907_ (.A1(_09418_),
    .A2(_09422_),
    .B1(_09546_),
    .C1(_09542_),
    .X(_09548_));
 sky130_fd_sc_hd__and2b_1 _16908_ (.A_N(_09547_),
    .B(_09548_),
    .X(_09549_));
 sky130_fd_sc_hd__xor2_2 _16909_ (.A(_09539_),
    .B(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__and2_1 _16910_ (.A(_08237_),
    .B(_09279_),
    .X(_09551_));
 sky130_fd_sc_hd__buf_2 _16911_ (.A(_09551_),
    .X(_09552_));
 sky130_fd_sc_hd__nor2_2 _16912_ (.A(_09117_),
    .B(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__inv_2 _16913_ (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_09554_));
 sky130_fd_sc_hd__mux2_2 _16914_ (.A0(_09554_),
    .A1(_09138_),
    .S(_05198_),
    .X(_09555_));
 sky130_fd_sc_hd__or3b_1 _16915_ (.A(_08873_),
    .B(_09555_),
    .C_N(_09421_),
    .X(_09556_));
 sky130_fd_sc_hd__o22ai_1 _16916_ (.A1(_08873_),
    .A2(_09540_),
    .B1(_09555_),
    .B2(_08872_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(_09556_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__xnor2_2 _16918_ (.A(_09553_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__or4_1 _16919_ (.A(_07602_),
    .B(_09283_),
    .C(_05209_),
    .D(_09287_),
    .X(_09560_));
 sky130_fd_sc_hd__or4_1 _16920_ (.A(_07598_),
    .B(_09283_),
    .C(_05210_),
    .D(_09433_),
    .X(_09561_));
 sky130_fd_sc_hd__xor2_1 _16921_ (.A(_09560_),
    .B(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__o31a_1 _16922_ (.A1(_07575_),
    .A2(_08983_),
    .A3(_09430_),
    .B1(_07586_),
    .X(_09563_));
 sky130_fd_sc_hd__a211o_1 _16923_ (.A1(_07585_),
    .A2(_09431_),
    .B1(_09563_),
    .C1(_09085_),
    .X(_09564_));
 sky130_fd_sc_hd__a22oi_4 _16924_ (.A1(_09283_),
    .A2(\rbzero.wall_tracer.stepDistY[10] ),
    .B1(_08235_),
    .B2(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__nor2_2 _16925_ (.A(_08816_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__xnor2_2 _16926_ (.A(_09562_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nor3_1 _16927_ (.A(_08215_),
    .B(_09294_),
    .C(_09427_),
    .Y(_09568_));
 sky130_fd_sc_hd__a21oi_2 _16928_ (.A1(_09428_),
    .A2(_09435_),
    .B1(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__xor2_2 _16929_ (.A(_09567_),
    .B(_09569_),
    .X(_09570_));
 sky130_fd_sc_hd__xnor2_2 _16930_ (.A(_09559_),
    .B(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__and2b_1 _16931_ (.A_N(_09436_),
    .B(_09437_),
    .X(_09572_));
 sky130_fd_sc_hd__a21o_1 _16932_ (.A1(_09425_),
    .A2(_09438_),
    .B1(_09572_),
    .X(_09573_));
 sky130_fd_sc_hd__xnor2_2 _16933_ (.A(_09571_),
    .B(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__xnor2_2 _16934_ (.A(_09550_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__nor2_1 _16935_ (.A(_09439_),
    .B(_09440_),
    .Y(_09576_));
 sky130_fd_sc_hd__a21o_1 _16936_ (.A1(_09415_),
    .A2(_09441_),
    .B1(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__xnor2_1 _16937_ (.A(_09575_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__xnor2_1 _16938_ (.A(_09538_),
    .B(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__nor2_1 _16939_ (.A(_09442_),
    .B(_09443_),
    .Y(_09580_));
 sky130_fd_sc_hd__a21o_1 _16940_ (.A1(_09405_),
    .A2(_09444_),
    .B1(_09580_),
    .X(_09581_));
 sky130_fd_sc_hd__xnor2_1 _16941_ (.A(_09579_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__xnor2_1 _16942_ (.A(_09517_),
    .B(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__nor2_1 _16943_ (.A(_09445_),
    .B(_09446_),
    .Y(_09584_));
 sky130_fd_sc_hd__a21oi_1 _16944_ (.A1(_09382_),
    .A2(_09447_),
    .B1(_09584_),
    .Y(_09585_));
 sky130_fd_sc_hd__xor2_1 _16945_ (.A(_09583_),
    .B(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__xnor2_1 _16946_ (.A(_09476_),
    .B(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__nor2_1 _16947_ (.A(_09448_),
    .B(_09449_),
    .Y(_09588_));
 sky130_fd_sc_hd__a21oi_1 _16948_ (.A1(_09347_),
    .A2(_09450_),
    .B1(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__xor2_1 _16949_ (.A(_09587_),
    .B(_09589_),
    .X(_09590_));
 sky130_fd_sc_hd__xor2_1 _16950_ (.A(_09345_),
    .B(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__and2_1 _16951_ (.A(_09454_),
    .B(_09591_),
    .X(_09592_));
 sky130_fd_sc_hd__nor2_1 _16952_ (.A(_09454_),
    .B(_09591_),
    .Y(_09593_));
 sky130_fd_sc_hd__nor2_4 _16953_ (.A(_09592_),
    .B(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__a21oi_1 _16954_ (.A1(_09342_),
    .A2(_09328_),
    .B1(_09456_),
    .Y(_09595_));
 sky130_fd_sc_hd__a31o_2 _16955_ (.A1(_09207_),
    .A2(_09330_),
    .A3(_09457_),
    .B1(_09595_),
    .X(_09596_));
 sky130_fd_sc_hd__xor2_4 _16956_ (.A(_09594_),
    .B(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__mux2_1 _16957_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_07895_),
    .X(_09598_));
 sky130_fd_sc_hd__nor2_1 _16958_ (.A(_09597_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__and2_1 _16959_ (.A(_09597_),
    .B(_09598_),
    .X(_09600_));
 sky130_fd_sc_hd__nor2_1 _16960_ (.A(_09599_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__xnor2_1 _16961_ (.A(_09082_),
    .B(_09601_),
    .Y(_09602_));
 sky130_fd_sc_hd__xnor2_1 _16962_ (.A(_09470_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__nand2_1 _16963_ (.A(_09085_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__o211a_1 _16964_ (.A1(\rbzero.wall_tracer.texu[4] ),
    .A2(_09085_),
    .B1(_04035_),
    .C1(_09604_),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_1 _16965_ (.A(_09587_),
    .B(_09589_),
    .Y(_09605_));
 sky130_fd_sc_hd__and2_1 _16966_ (.A(_09345_),
    .B(_09590_),
    .X(_09606_));
 sky130_fd_sc_hd__or2b_1 _16967_ (.A(_09516_),
    .B_N(_09477_),
    .X(_09607_));
 sky130_fd_sc_hd__xnor2_1 _16968_ (.A(_09486_),
    .B(_09495_),
    .Y(_09608_));
 sky130_fd_sc_hd__a31o_1 _16969_ (.A1(_09485_),
    .A2(_09486_),
    .A3(_09497_),
    .B1(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(\rbzero.wall_tracer.visualWallDist[11] ),
    .B(_04015_),
    .Y(_09610_));
 sky130_fd_sc_hd__nor2_2 _16971_ (.A(_05211_),
    .B(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__and2_1 _16972_ (.A(_08162_),
    .B(_09611_),
    .X(_09612_));
 sky130_fd_sc_hd__xnor2_2 _16973_ (.A(_09609_),
    .B(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__a21oi_4 _16974_ (.A1(_09514_),
    .A2(_09607_),
    .B1(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__and3_1 _16975_ (.A(_09514_),
    .B(_09607_),
    .C(_09613_),
    .X(_09615_));
 sky130_fd_sc_hd__nor2_1 _16976_ (.A(_09614_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__a21o_1 _16977_ (.A1(_09498_),
    .A2(_09512_),
    .B1(_09510_),
    .X(_09617_));
 sky130_fd_sc_hd__or2b_1 _16978_ (.A(_09536_),
    .B_N(_09520_),
    .X(_09618_));
 sky130_fd_sc_hd__or2b_1 _16979_ (.A(_09537_),
    .B_N(_09518_),
    .X(_09619_));
 sky130_fd_sc_hd__nor2_1 _16980_ (.A(_08160_),
    .B(_09483_),
    .Y(_09620_));
 sky130_fd_sc_hd__nor2_1 _16981_ (.A(_05211_),
    .B(_09350_),
    .Y(_09621_));
 sky130_fd_sc_hd__o22a_1 _16982_ (.A1(_08329_),
    .A2(_09216_),
    .B1(_09351_),
    .B2(_08054_),
    .X(_09622_));
 sky130_fd_sc_hd__a31oi_1 _16983_ (.A1(_08331_),
    .A2(_09621_),
    .A3(_09488_),
    .B1(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(_09620_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__or2_1 _16985_ (.A(_09620_),
    .B(_09623_),
    .X(_09625_));
 sky130_fd_sc_hd__and2_1 _16986_ (.A(_09624_),
    .B(_09625_),
    .X(_09626_));
 sky130_fd_sc_hd__nor2_1 _16987_ (.A(_08823_),
    .B(_09164_),
    .Y(_09627_));
 sky130_fd_sc_hd__o22a_1 _16988_ (.A1(_08821_),
    .A2(_09028_),
    .B1(_08425_),
    .B2(_09243_),
    .X(_09628_));
 sky130_fd_sc_hd__or4_1 _16989_ (.A(_08075_),
    .B(_08821_),
    .C(_09028_),
    .D(_08425_),
    .X(_09629_));
 sky130_fd_sc_hd__and2b_1 _16990_ (.A_N(_09628_),
    .B(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__xnor2_1 _16991_ (.A(_09627_),
    .B(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__o31a_1 _16992_ (.A1(_08335_),
    .A2(_09217_),
    .A3(_09489_),
    .B1(_09490_),
    .X(_09632_));
 sky130_fd_sc_hd__or2_1 _16993_ (.A(_09631_),
    .B(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__nand2_1 _16994_ (.A(_09631_),
    .B(_09632_),
    .Y(_09634_));
 sky130_fd_sc_hd__and2_1 _16995_ (.A(_09633_),
    .B(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__nand2_1 _16996_ (.A(_09626_),
    .B(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__or2_1 _16997_ (.A(_09626_),
    .B(_09635_),
    .X(_09637_));
 sky130_fd_sc_hd__and2_1 _16998_ (.A(_09636_),
    .B(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__a21bo_1 _16999_ (.A1(_09501_),
    .A2(_09504_),
    .B1_N(_09503_),
    .X(_09639_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_09521_),
    .B(_09525_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _17001_ (.A(_09245_),
    .B(_08159_),
    .Y(_09641_));
 sky130_fd_sc_hd__o22a_1 _17002_ (.A1(_07994_),
    .A2(_08058_),
    .B1(_08151_),
    .B2(_08705_),
    .X(_09642_));
 sky130_fd_sc_hd__or4_1 _17003_ (.A(_07994_),
    .B(_08705_),
    .C(_08058_),
    .D(_08150_),
    .X(_09643_));
 sky130_fd_sc_hd__and2b_1 _17004_ (.A_N(_09642_),
    .B(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__xnor2_1 _17005_ (.A(_09641_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__xnor2_1 _17006_ (.A(_09640_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__xnor2_1 _17007_ (.A(_09639_),
    .B(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__a21oi_1 _17008_ (.A1(_09387_),
    .A2(_09390_),
    .B1(_09505_),
    .Y(_09648_));
 sky130_fd_sc_hd__a21oi_1 _17009_ (.A1(_09499_),
    .A2(_09506_),
    .B1(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__nor2_1 _17010_ (.A(_09647_),
    .B(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__and2_1 _17011_ (.A(_09647_),
    .B(_09649_),
    .X(_09651_));
 sky130_fd_sc_hd__nor2_1 _17012_ (.A(_09650_),
    .B(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__xnor2_1 _17013_ (.A(_09638_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__a21o_1 _17014_ (.A1(_09618_),
    .A2(_09619_),
    .B1(_09653_),
    .X(_09654_));
 sky130_fd_sc_hd__nand3_1 _17015_ (.A(_09618_),
    .B(_09619_),
    .C(_09653_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _17016_ (.A(_09654_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__xnor2_2 _17017_ (.A(_09617_),
    .B(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__nor2_1 _17018_ (.A(_09533_),
    .B(_09534_),
    .Y(_09658_));
 sky130_fd_sc_hd__a21o_1 _17019_ (.A1(_09528_),
    .A2(_09535_),
    .B1(_09658_),
    .X(_09659_));
 sky130_fd_sc_hd__a21o_2 _17020_ (.A1(_09539_),
    .A2(_09548_),
    .B1(_09547_),
    .X(_09660_));
 sky130_fd_sc_hd__clkbuf_4 _17021_ (.A(_07976_),
    .X(_09661_));
 sky130_fd_sc_hd__o22ai_1 _17022_ (.A1(_08204_),
    .A2(_09103_),
    .B1(_08493_),
    .B2(_08383_),
    .Y(_09662_));
 sky130_fd_sc_hd__a21o_1 _17023_ (.A1(_08202_),
    .A2(_08203_),
    .B1(_08129_),
    .X(_09663_));
 sky130_fd_sc_hd__or3_1 _17024_ (.A(_08383_),
    .B(_09103_),
    .C(_09663_),
    .X(_09664_));
 sky130_fd_sc_hd__or4bb_2 _17025_ (.A(_09661_),
    .B(_08047_),
    .C_N(_09662_),
    .D_N(_09664_),
    .X(_09665_));
 sky130_fd_sc_hd__a2bb2o_1 _17026_ (.A1_N(_09661_),
    .A2_N(_08047_),
    .B1(_09662_),
    .B2(_09664_),
    .X(_09666_));
 sky130_fd_sc_hd__nand2_1 _17027_ (.A(_09665_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__buf_4 _17028_ (.A(_08570_),
    .X(_09668_));
 sky130_fd_sc_hd__nor2_2 _17029_ (.A(_08178_),
    .B(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__nor2_4 _17030_ (.A(_09276_),
    .B(_08111_),
    .Y(_09670_));
 sky130_fd_sc_hd__o22a_1 _17031_ (.A1(_07959_),
    .A2(_09276_),
    .B1(_08111_),
    .B2(_09126_),
    .X(_09671_));
 sky130_fd_sc_hd__a21oi_2 _17032_ (.A1(_09545_),
    .A2(_09670_),
    .B1(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__xnor2_2 _17033_ (.A(_09669_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__clkbuf_4 _17034_ (.A(_09103_),
    .X(_09674_));
 sky130_fd_sc_hd__nand2_1 _17035_ (.A(_09396_),
    .B(_09669_),
    .Y(_09675_));
 sky130_fd_sc_hd__o31a_1 _17036_ (.A1(_08383_),
    .A2(_09674_),
    .A3(_09531_),
    .B1(_09675_),
    .X(_09676_));
 sky130_fd_sc_hd__xor2_2 _17037_ (.A(_09673_),
    .B(_09676_),
    .X(_09677_));
 sky130_fd_sc_hd__xor2_2 _17038_ (.A(_09667_),
    .B(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__xor2_2 _17039_ (.A(_09660_),
    .B(_09678_),
    .X(_09679_));
 sky130_fd_sc_hd__xnor2_2 _17040_ (.A(_09659_),
    .B(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__or3_1 _17041_ (.A(_09114_),
    .B(_09126_),
    .C(_09544_),
    .X(_09681_));
 sky130_fd_sc_hd__a21bo_2 _17042_ (.A1(_09409_),
    .A2(_09543_),
    .B1_N(_09681_),
    .X(_09682_));
 sky130_fd_sc_hd__a21bo_1 _17043_ (.A1(_09553_),
    .A2(_09557_),
    .B1_N(_09556_),
    .X(_09683_));
 sky130_fd_sc_hd__nor2_1 _17044_ (.A(_08767_),
    .B(_09417_),
    .Y(_09684_));
 sky130_fd_sc_hd__a21o_1 _17045_ (.A1(_09141_),
    .A2(_09420_),
    .B1(_08194_),
    .X(_09685_));
 sky130_fd_sc_hd__a21oi_2 _17046_ (.A1(_08237_),
    .A2(_09279_),
    .B1(_08283_),
    .Y(_09686_));
 sky130_fd_sc_hd__xnor2_1 _17047_ (.A(_09685_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__xor2_1 _17048_ (.A(_09684_),
    .B(_09687_),
    .X(_09688_));
 sky130_fd_sc_hd__and2_1 _17049_ (.A(_09683_),
    .B(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__or2_1 _17050_ (.A(_09683_),
    .B(_09688_),
    .X(_09690_));
 sky130_fd_sc_hd__or2b_1 _17051_ (.A(_09689_),
    .B_N(_09690_),
    .X(_09691_));
 sky130_fd_sc_hd__xnor2_4 _17052_ (.A(_09682_),
    .B(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__buf_4 _17053_ (.A(_09555_),
    .X(_09693_));
 sky130_fd_sc_hd__nor2_2 _17054_ (.A(_08873_),
    .B(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__nand2_4 _17055_ (.A(_05210_),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_09695_));
 sky130_fd_sc_hd__a21oi_2 _17056_ (.A1(_09292_),
    .A2(_09695_),
    .B1(_08872_),
    .Y(_09696_));
 sky130_fd_sc_hd__inv_2 _17057_ (.A(_07589_),
    .Y(_09697_));
 sky130_fd_sc_hd__a31o_1 _17058_ (.A1(_07585_),
    .A2(_09697_),
    .A3(_09431_),
    .B1(_09085_),
    .X(_09698_));
 sky130_fd_sc_hd__a22oi_4 _17059_ (.A1(_09283_),
    .A2(\rbzero.wall_tracer.stepDistY[11] ),
    .B1(_08235_),
    .B2(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__or2_2 _17060_ (.A(_08816_),
    .B(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__xnor2_2 _17061_ (.A(_09696_),
    .B(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__xor2_4 _17062_ (.A(_09694_),
    .B(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__nor2_4 _17063_ (.A(_03953_),
    .B(_09283_),
    .Y(_09703_));
 sky130_fd_sc_hd__nand2_4 _17064_ (.A(_05198_),
    .B(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__or4_1 _17065_ (.A(_07602_),
    .B(_09283_),
    .C(_05210_),
    .D(_09433_),
    .X(_09705_));
 sky130_fd_sc_hd__or4_1 _17066_ (.A(_03953_),
    .B(_09283_),
    .C(_08377_),
    .D(_09433_),
    .X(_09706_));
 sky130_fd_sc_hd__a21bo_2 _17067_ (.A1(_09704_),
    .A2(_09705_),
    .B1_N(_09706_),
    .X(_09707_));
 sky130_fd_sc_hd__or2_2 _17068_ (.A(_08519_),
    .B(_09565_),
    .X(_09708_));
 sky130_fd_sc_hd__xnor2_4 _17069_ (.A(_09707_),
    .B(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(_09560_),
    .B(_09561_),
    .Y(_09710_));
 sky130_fd_sc_hd__nor2_1 _17071_ (.A(_09560_),
    .B(_09561_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21oi_4 _17072_ (.A1(_09710_),
    .A2(_09566_),
    .B1(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__xor2_4 _17073_ (.A(_09709_),
    .B(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__xnor2_4 _17074_ (.A(_09702_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__nor2_1 _17075_ (.A(_09567_),
    .B(_09569_),
    .Y(_09715_));
 sky130_fd_sc_hd__a21oi_2 _17076_ (.A1(_09559_),
    .A2(_09570_),
    .B1(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__xor2_4 _17077_ (.A(_09714_),
    .B(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__xnor2_4 _17078_ (.A(_09692_),
    .B(_09717_),
    .Y(_09718_));
 sky130_fd_sc_hd__and2b_1 _17079_ (.A_N(_09571_),
    .B(_09573_),
    .X(_09719_));
 sky130_fd_sc_hd__a21oi_2 _17080_ (.A1(_09550_),
    .A2(_09574_),
    .B1(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__xor2_4 _17081_ (.A(_09718_),
    .B(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__xnor2_2 _17082_ (.A(_09680_),
    .B(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__or2b_1 _17083_ (.A(_09575_),
    .B_N(_09577_),
    .X(_09723_));
 sky130_fd_sc_hd__a21boi_2 _17084_ (.A1(_09538_),
    .A2(_09578_),
    .B1_N(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__xor2_2 _17085_ (.A(_09722_),
    .B(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__xnor2_2 _17086_ (.A(_09657_),
    .B(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__and2b_1 _17087_ (.A_N(_09579_),
    .B(_09581_),
    .X(_09727_));
 sky130_fd_sc_hd__a21oi_2 _17088_ (.A1(_09517_),
    .A2(_09582_),
    .B1(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__xor2_2 _17089_ (.A(_09726_),
    .B(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__xnor2_2 _17090_ (.A(_09616_),
    .B(_09729_),
    .Y(_09730_));
 sky130_fd_sc_hd__nor2_1 _17091_ (.A(_09583_),
    .B(_09585_),
    .Y(_09731_));
 sky130_fd_sc_hd__a21oi_2 _17092_ (.A1(_09476_),
    .A2(_09586_),
    .B1(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__xor2_2 _17093_ (.A(_09730_),
    .B(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__xor2_1 _17094_ (.A(_09474_),
    .B(_09733_),
    .X(_09734_));
 sky130_fd_sc_hd__nor3_1 _17095_ (.A(_09605_),
    .B(_09606_),
    .C(_09734_),
    .Y(_09735_));
 sky130_fd_sc_hd__o21a_1 _17096_ (.A1(_09605_),
    .A2(_09606_),
    .B1(_09734_),
    .X(_09736_));
 sky130_fd_sc_hd__nor2_2 _17097_ (.A(_09735_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__a21oi_2 _17098_ (.A1(_09594_),
    .A2(_09596_),
    .B1(_09592_),
    .Y(_09738_));
 sky130_fd_sc_hd__xnor2_4 _17099_ (.A(_09737_),
    .B(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__mux2_1 _17100_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_07895_),
    .X(_09740_));
 sky130_fd_sc_hd__xnor2_2 _17101_ (.A(_09082_),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__xnor2_1 _17102_ (.A(_09739_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__inv_2 _17103_ (.A(_09599_),
    .Y(_09743_));
 sky130_fd_sc_hd__o311a_1 _17104_ (.A1(_09461_),
    .A2(_09465_),
    .A3(_09600_),
    .B1(_09742_),
    .C1(_09743_),
    .X(_09744_));
 sky130_fd_sc_hd__a211o_1 _17105_ (.A1(_09470_),
    .A2(_09743_),
    .B1(_09600_),
    .C1(_09742_),
    .X(_09745_));
 sky130_fd_sc_hd__or3b_1 _17106_ (.A(_05194_),
    .B(_09744_),
    .C_N(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__o211a_1 _17107_ (.A1(\rbzero.wall_tracer.texu[5] ),
    .A2(_09085_),
    .B1(_04035_),
    .C1(_09746_),
    .X(_00516_));
 sky130_fd_sc_hd__or2_1 _17108_ (.A(_03555_),
    .B(_04037_),
    .X(_09747_));
 sky130_fd_sc_hd__clkbuf_2 _17109_ (.A(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__nor2_1 _17110_ (.A(_03474_),
    .B(_09748_),
    .Y(_00517_));
 sky130_fd_sc_hd__nor2_1 _17111_ (.A(_03555_),
    .B(_04037_),
    .Y(_09749_));
 sky130_fd_sc_hd__clkbuf_4 _17112_ (.A(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__or2_1 _17113_ (.A(_04814_),
    .B(_03474_),
    .X(_09751_));
 sky130_fd_sc_hd__and3_1 _17114_ (.A(_04821_),
    .B(_09750_),
    .C(_09751_),
    .X(_09752_));
 sky130_fd_sc_hd__clkbuf_1 _17115_ (.A(_09752_),
    .X(_00518_));
 sky130_fd_sc_hd__buf_6 _17116_ (.A(_05189_),
    .X(_09753_));
 sky130_fd_sc_hd__a21o_1 _17117_ (.A1(_04814_),
    .A2(_03474_),
    .B1(_04317_),
    .X(_09754_));
 sky130_fd_sc_hd__and3_1 _17118_ (.A(_09753_),
    .B(_04319_),
    .C(_09754_),
    .X(_09755_));
 sky130_fd_sc_hd__clkbuf_1 _17119_ (.A(_09755_),
    .X(_00519_));
 sky130_fd_sc_hd__nor2_1 _17120_ (.A(_04417_),
    .B(_09748_),
    .Y(_00520_));
 sky130_fd_sc_hd__nor2_1 _17121_ (.A(_04426_),
    .B(_09748_),
    .Y(_00521_));
 sky130_fd_sc_hd__and2_1 _17122_ (.A(_04430_),
    .B(_09750_),
    .X(_09756_));
 sky130_fd_sc_hd__clkbuf_1 _17123_ (.A(_09756_),
    .X(_00522_));
 sky130_fd_sc_hd__nor2_1 _17124_ (.A(_04422_),
    .B(_09748_),
    .Y(_00523_));
 sky130_fd_sc_hd__and2_1 _17125_ (.A(_04443_),
    .B(_09750_),
    .X(_09757_));
 sky130_fd_sc_hd__clkbuf_1 _17126_ (.A(_09757_),
    .X(_00524_));
 sky130_fd_sc_hd__or2_1 _17127_ (.A(_04154_),
    .B(_04442_),
    .X(_09758_));
 sky130_fd_sc_hd__and3_1 _17128_ (.A(_04446_),
    .B(_09750_),
    .C(_09758_),
    .X(_09759_));
 sky130_fd_sc_hd__clkbuf_1 _17129_ (.A(_09759_),
    .X(_00525_));
 sky130_fd_sc_hd__or2_1 _17130_ (.A(_03477_),
    .B(_04446_),
    .X(_09760_));
 sky130_fd_sc_hd__nand2_1 _17131_ (.A(_03477_),
    .B(_04446_),
    .Y(_09761_));
 sky130_fd_sc_hd__a21oi_1 _17132_ (.A1(_09760_),
    .A2(_09761_),
    .B1(_09748_),
    .Y(_00526_));
 sky130_fd_sc_hd__clkbuf_8 _17133_ (.A(_07706_),
    .X(_09762_));
 sky130_fd_sc_hd__a22o_1 _17134_ (.A1(\rbzero.row_render.side ),
    .A2(_09762_),
    .B1(_07728_),
    .B2(_07895_),
    .X(_00527_));
 sky130_fd_sc_hd__buf_2 _17135_ (.A(_07831_),
    .X(_09763_));
 sky130_fd_sc_hd__buf_2 _17136_ (.A(_07855_),
    .X(_09764_));
 sky130_fd_sc_hd__a2bb2o_1 _17137_ (.A1_N(_07514_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[0] ),
    .B2(_09764_),
    .X(_00528_));
 sky130_fd_sc_hd__a2bb2o_1 _17138_ (.A1_N(_07524_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[1] ),
    .B2(_09764_),
    .X(_00529_));
 sky130_fd_sc_hd__a2bb2o_1 _17139_ (.A1_N(_07530_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[2] ),
    .B2(_09764_),
    .X(_00530_));
 sky130_fd_sc_hd__a2bb2o_1 _17140_ (.A1_N(_07536_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[3] ),
    .B2(_09764_),
    .X(_00531_));
 sky130_fd_sc_hd__a22o_1 _17141_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_09762_),
    .B1(_07541_),
    .B2(_07756_),
    .X(_00532_));
 sky130_fd_sc_hd__nor2_2 _17142_ (.A(_07468_),
    .B(_07544_),
    .Y(_09765_));
 sky130_fd_sc_hd__a2bb2o_1 _17143_ (.A1_N(_09765_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[5] ),
    .B2(_09764_),
    .X(_00533_));
 sky130_fd_sc_hd__a2bb2o_1 _17144_ (.A1_N(_07549_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[6] ),
    .B2(_09764_),
    .X(_00534_));
 sky130_fd_sc_hd__a2bb2o_1 _17145_ (.A1_N(_07552_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[7] ),
    .B2(_09764_),
    .X(_00535_));
 sky130_fd_sc_hd__a2bb2o_1 _17146_ (.A1_N(_07555_),
    .A2_N(_09763_),
    .B1(\rbzero.row_render.size[8] ),
    .B2(_09764_),
    .X(_00536_));
 sky130_fd_sc_hd__a22o_1 _17147_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_09762_),
    .B1(_07560_),
    .B2(_07756_),
    .X(_00537_));
 sky130_fd_sc_hd__a22o_1 _17148_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_09762_),
    .B1(_07562_),
    .B2(_07756_),
    .X(_00538_));
 sky130_fd_sc_hd__a22o_1 _17149_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_09762_),
    .B1(_07728_),
    .B2(\rbzero.wall_tracer.texu[0] ),
    .X(_00539_));
 sky130_fd_sc_hd__buf_4 _17150_ (.A(_07706_),
    .X(_09766_));
 sky130_fd_sc_hd__a22o_1 _17151_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_09766_),
    .B1(_07728_),
    .B2(\rbzero.wall_tracer.texu[1] ),
    .X(_00540_));
 sky130_fd_sc_hd__a22o_1 _17152_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_09766_),
    .B1(_07728_),
    .B2(\rbzero.wall_tracer.texu[2] ),
    .X(_00541_));
 sky130_fd_sc_hd__a22o_1 _17153_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_09766_),
    .B1(_07728_),
    .B2(net511),
    .X(_00542_));
 sky130_fd_sc_hd__a22o_1 _17154_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_09766_),
    .B1(_07728_),
    .B2(\rbzero.wall_tracer.texu[4] ),
    .X(_00543_));
 sky130_fd_sc_hd__a22o_1 _17155_ (.A1(\rbzero.row_render.texu[5] ),
    .A2(_09766_),
    .B1(_07728_),
    .B2(\rbzero.wall_tracer.texu[5] ),
    .X(_00544_));
 sky130_fd_sc_hd__clkbuf_4 _17156_ (.A(_07679_),
    .X(_09767_));
 sky130_fd_sc_hd__a22o_1 _17157_ (.A1(\rbzero.traced_texa[-12] ),
    .A2(_09766_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-12] ),
    .X(_00545_));
 sky130_fd_sc_hd__a22o_1 _17158_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_09766_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00546_));
 sky130_fd_sc_hd__a22o_1 _17159_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_09766_),
    .B1(_09767_),
    .B2(_07601_),
    .X(_00547_));
 sky130_fd_sc_hd__a22o_1 _17160_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_09766_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00548_));
 sky130_fd_sc_hd__a22o_1 _17161_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_09766_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00549_));
 sky130_fd_sc_hd__clkbuf_4 _17162_ (.A(_07706_),
    .X(_09768_));
 sky130_fd_sc_hd__a22o_1 _17163_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_09768_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00550_));
 sky130_fd_sc_hd__a22o_1 _17164_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_09768_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00551_));
 sky130_fd_sc_hd__a22o_1 _17165_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_09768_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00552_));
 sky130_fd_sc_hd__a22o_1 _17166_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_09768_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00553_));
 sky130_fd_sc_hd__a22o_1 _17167_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_09768_),
    .B1(_09767_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00554_));
 sky130_fd_sc_hd__clkbuf_4 _17168_ (.A(_07679_),
    .X(_09769_));
 sky130_fd_sc_hd__a22o_1 _17169_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_09768_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00555_));
 sky130_fd_sc_hd__a22o_1 _17170_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_09768_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00556_));
 sky130_fd_sc_hd__a22o_1 _17171_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_09768_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00557_));
 sky130_fd_sc_hd__a22o_1 _17172_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_09768_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00558_));
 sky130_fd_sc_hd__a22o_1 _17173_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_09768_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00559_));
 sky130_fd_sc_hd__clkbuf_4 _17174_ (.A(_07706_),
    .X(_09770_));
 sky130_fd_sc_hd__a22o_1 _17175_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_09770_),
    .B1(_09769_),
    .B2(net514),
    .X(_00560_));
 sky130_fd_sc_hd__a22o_1 _17176_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_09770_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00561_));
 sky130_fd_sc_hd__a22o_1 _17177_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_09770_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00562_));
 sky130_fd_sc_hd__a22o_1 _17178_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_09770_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00563_));
 sky130_fd_sc_hd__a22o_1 _17179_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_09770_),
    .B1(_09769_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00564_));
 sky130_fd_sc_hd__clkbuf_4 _17180_ (.A(_07679_),
    .X(_09771_));
 sky130_fd_sc_hd__a22o_1 _17181_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_09770_),
    .B1(_09771_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00565_));
 sky130_fd_sc_hd__a22o_1 _17182_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_09770_),
    .B1(_09771_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00566_));
 sky130_fd_sc_hd__a22o_1 _17183_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_09770_),
    .B1(_09771_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00567_));
 sky130_fd_sc_hd__a22o_1 _17184_ (.A1(\rbzero.traced_texa[11] ),
    .A2(_09770_),
    .B1(_09771_),
    .B2(\rbzero.wall_tracer.visualWallDist[11] ),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _17185_ (.A0(\rbzero.wall_tracer.wall[0] ),
    .A1(\rbzero.row_render.wall[0] ),
    .S(_07830_),
    .X(_09772_));
 sky130_fd_sc_hd__clkbuf_1 _17186_ (.A(_09772_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(\rbzero.wall_tracer.wall[1] ),
    .A1(\rbzero.row_render.wall[1] ),
    .S(_07830_),
    .X(_09773_));
 sky130_fd_sc_hd__clkbuf_1 _17188_ (.A(_09773_),
    .X(_00570_));
 sky130_fd_sc_hd__xor2_1 _17189_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_05512_),
    .X(_09774_));
 sky130_fd_sc_hd__a21o_1 _17190_ (.A1(\rbzero.wall_tracer.mapX[5] ),
    .A2(_05512_),
    .B1(_05527_),
    .X(_09775_));
 sky130_fd_sc_hd__o21a_1 _17191_ (.A1(\rbzero.wall_tracer.mapX[5] ),
    .A2(_05512_),
    .B1(_09775_),
    .X(_09776_));
 sky130_fd_sc_hd__or2_1 _17192_ (.A(_09774_),
    .B(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__nand2_1 _17193_ (.A(_09774_),
    .B(_09776_),
    .Y(_09778_));
 sky130_fd_sc_hd__nor2_4 _17194_ (.A(_04019_),
    .B(_05412_),
    .Y(_09779_));
 sky130_fd_sc_hd__inv_2 _17195_ (.A(_05413_),
    .Y(_09780_));
 sky130_fd_sc_hd__buf_6 _17196_ (.A(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__a32o_1 _17197_ (.A1(_09777_),
    .A2(_09778_),
    .A3(_09779_),
    .B1(_09781_),
    .B2(\rbzero.wall_tracer.mapX[6] ),
    .X(_00571_));
 sky130_fd_sc_hd__a21bo_1 _17198_ (.A1(\rbzero.wall_tracer.mapX[6] ),
    .A2(_05512_),
    .B1_N(_09778_),
    .X(_09782_));
 sky130_fd_sc_hd__and2_1 _17199_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_05512_),
    .X(_09783_));
 sky130_fd_sc_hd__nor2_1 _17200_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_05525_),
    .Y(_09784_));
 sky130_fd_sc_hd__or2_1 _17201_ (.A(_09783_),
    .B(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__xnor2_1 _17202_ (.A(_09782_),
    .B(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__a22o_1 _17203_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(_09781_),
    .B1(_09779_),
    .B2(_09786_),
    .X(_00572_));
 sky130_fd_sc_hd__o21a_1 _17204_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(_05512_),
    .B1(_09782_),
    .X(_09787_));
 sky130_fd_sc_hd__xor2_1 _17205_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_05525_),
    .X(_09788_));
 sky130_fd_sc_hd__or3_1 _17206_ (.A(_09783_),
    .B(_09787_),
    .C(_09788_),
    .X(_09789_));
 sky130_fd_sc_hd__o21ai_1 _17207_ (.A1(_09783_),
    .A2(_09787_),
    .B1(_09788_),
    .Y(_09790_));
 sky130_fd_sc_hd__a32o_1 _17208_ (.A1(_09779_),
    .A2(_09789_),
    .A3(_09790_),
    .B1(_09781_),
    .B2(\rbzero.wall_tracer.mapX[8] ),
    .X(_00573_));
 sky130_fd_sc_hd__a21bo_1 _17209_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_05525_),
    .B1_N(_09790_),
    .X(_09791_));
 sky130_fd_sc_hd__and2_1 _17210_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_05525_),
    .X(_09792_));
 sky130_fd_sc_hd__nor2_1 _17211_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_05525_),
    .Y(_09793_));
 sky130_fd_sc_hd__or2_1 _17212_ (.A(_09792_),
    .B(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__xnor2_1 _17213_ (.A(_09791_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__a22o_1 _17214_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09781_),
    .B1(_09779_),
    .B2(_09795_),
    .X(_00574_));
 sky130_fd_sc_hd__o21a_1 _17215_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_05525_),
    .B1(_09791_),
    .X(_09796_));
 sky130_fd_sc_hd__xor2_1 _17216_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(_05525_),
    .X(_09797_));
 sky130_fd_sc_hd__or3_1 _17217_ (.A(_09792_),
    .B(_09796_),
    .C(_09797_),
    .X(_09798_));
 sky130_fd_sc_hd__o21ai_1 _17218_ (.A1(_09792_),
    .A2(_09796_),
    .B1(_09797_),
    .Y(_09799_));
 sky130_fd_sc_hd__a32o_1 _17219_ (.A1(_09779_),
    .A2(_09798_),
    .A3(_09799_),
    .B1(_09781_),
    .B2(\rbzero.wall_tracer.mapX[10] ),
    .X(_00575_));
 sky130_fd_sc_hd__a21bo_1 _17220_ (.A1(\rbzero.wall_tracer.mapX[10] ),
    .A2(_05525_),
    .B1_N(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__xnor2_1 _17221_ (.A(\rbzero.wall_tracer.mapX[11] ),
    .B(_05525_),
    .Y(_09801_));
 sky130_fd_sc_hd__xnor2_1 _17222_ (.A(_09800_),
    .B(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__a22o_1 _17223_ (.A1(\rbzero.wall_tracer.mapX[11] ),
    .A2(_09781_),
    .B1(_09779_),
    .B2(_09802_),
    .X(_00576_));
 sky130_fd_sc_hd__and2_1 _17224_ (.A(_08939_),
    .B(_08851_),
    .X(_09803_));
 sky130_fd_sc_hd__xor2_1 _17225_ (.A(_08937_),
    .B(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__and3_1 _17226_ (.A(_08939_),
    .B(_08850_),
    .C(_08936_),
    .X(_09805_));
 sky130_fd_sc_hd__nor2_1 _17227_ (.A(_09804_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__buf_6 _17228_ (.A(_05203_),
    .X(_09807_));
 sky130_fd_sc_hd__a211o_1 _17229_ (.A1(_09804_),
    .A2(_09805_),
    .B1(_09806_),
    .C1(_09807_),
    .X(_09808_));
 sky130_fd_sc_hd__o21ai_1 _17230_ (.A1(\rbzero.wall_tracer.trackDistX[-12] ),
    .A2(\rbzero.wall_tracer.stepDistX[-12] ),
    .B1(_09807_),
    .Y(_09809_));
 sky130_fd_sc_hd__a21o_1 _17231_ (.A1(\rbzero.wall_tracer.trackDistX[-12] ),
    .A2(\rbzero.wall_tracer.stepDistX[-12] ),
    .B1(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__and3_1 _17232_ (.A(_05413_),
    .B(_09808_),
    .C(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__a21oi_1 _17233_ (.A1(_05243_),
    .A2(_09781_),
    .B1(_09811_),
    .Y(_00577_));
 sky130_fd_sc_hd__buf_4 _17234_ (.A(_04016_),
    .X(_09812_));
 sky130_fd_sc_hd__or2_1 _17235_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .X(_09813_));
 sky130_fd_sc_hd__nand2_1 _17236_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .Y(_09814_));
 sky130_fd_sc_hd__and4_1 _17237_ (.A(\rbzero.wall_tracer.trackDistX[-12] ),
    .B(\rbzero.wall_tracer.stepDistX[-12] ),
    .C(_09813_),
    .D(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__a22oi_1 _17238_ (.A1(\rbzero.wall_tracer.trackDistX[-12] ),
    .A2(\rbzero.wall_tracer.stepDistX[-12] ),
    .B1(_09813_),
    .B2(_09814_),
    .Y(_09816_));
 sky130_fd_sc_hd__buf_4 _17239_ (.A(_05413_),
    .X(_09817_));
 sky130_fd_sc_hd__a21oi_1 _17240_ (.A1(_08940_),
    .A2(_08943_),
    .B1(_05204_),
    .Y(_09818_));
 sky130_fd_sc_hd__o21ai_1 _17241_ (.A1(_08940_),
    .A2(_08943_),
    .B1(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__o311a_1 _17242_ (.A1(_09812_),
    .A2(_09815_),
    .A3(_09816_),
    .B1(_09817_),
    .C1(_09819_),
    .X(_09820_));
 sky130_fd_sc_hd__a21oi_1 _17243_ (.A1(_05242_),
    .A2(_09781_),
    .B1(_09820_),
    .Y(_00578_));
 sky130_fd_sc_hd__or2_1 _17244_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_09821_));
 sky130_fd_sc_hd__nand2_1 _17245_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_09822_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09815_),
    .X(_09823_));
 sky130_fd_sc_hd__a21oi_1 _17247_ (.A1(_09821_),
    .A2(_09822_),
    .B1(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__a31o_1 _17248_ (.A1(_09823_),
    .A2(_09821_),
    .A3(_09822_),
    .B1(_05531_),
    .X(_09825_));
 sky130_fd_sc_hd__o21ai_1 _17249_ (.A1(_08944_),
    .A2(_08948_),
    .B1(_04016_),
    .Y(_09826_));
 sky130_fd_sc_hd__a21o_1 _17250_ (.A1(_08944_),
    .A2(_08948_),
    .B1(_09826_),
    .X(_09827_));
 sky130_fd_sc_hd__o21ai_1 _17251_ (.A1(_09824_),
    .A2(_09825_),
    .B1(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__mux2_1 _17252_ (.A0(\rbzero.wall_tracer.trackDistX[-10] ),
    .A1(_09828_),
    .S(_05414_),
    .X(_09829_));
 sky130_fd_sc_hd__clkbuf_1 _17253_ (.A(_09829_),
    .X(_00579_));
 sky130_fd_sc_hd__or2_1 _17254_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_09830_));
 sky130_fd_sc_hd__nand2_1 _17255_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_09831_));
 sky130_fd_sc_hd__a21bo_1 _17256_ (.A1(_09823_),
    .A2(_09821_),
    .B1_N(_09822_),
    .X(_09832_));
 sky130_fd_sc_hd__and3_1 _17257_ (.A(_09830_),
    .B(_09831_),
    .C(_09832_),
    .X(_09833_));
 sky130_fd_sc_hd__a21oi_1 _17258_ (.A1(_09830_),
    .A2(_09831_),
    .B1(_09832_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_1 _17259_ (.A(_05531_),
    .B(_09069_),
    .Y(_09835_));
 sky130_fd_sc_hd__o31ai_1 _17260_ (.A1(_09812_),
    .A2(_09833_),
    .A3(_09834_),
    .B1(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__mux2_1 _17261_ (.A0(\rbzero.wall_tracer.trackDistX[-9] ),
    .A1(_09836_),
    .S(_05414_),
    .X(_09837_));
 sky130_fd_sc_hd__clkbuf_1 _17262_ (.A(_09837_),
    .X(_00580_));
 sky130_fd_sc_hd__nor2_1 _17263_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_09838_));
 sky130_fd_sc_hd__and2_1 _17264_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_09839_));
 sky130_fd_sc_hd__a21boi_1 _17265_ (.A1(_09830_),
    .A2(_09832_),
    .B1_N(_09831_),
    .Y(_09840_));
 sky130_fd_sc_hd__nor3_1 _17266_ (.A(_09838_),
    .B(_09839_),
    .C(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__o21a_1 _17267_ (.A1(_09838_),
    .A2(_09839_),
    .B1(_09840_),
    .X(_09842_));
 sky130_fd_sc_hd__nand2_1 _17268_ (.A(_05531_),
    .B(_09068_),
    .Y(_09843_));
 sky130_fd_sc_hd__o31ai_1 _17269_ (.A1(_09812_),
    .A2(_09841_),
    .A3(_09842_),
    .B1(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__mux2_1 _17270_ (.A0(\rbzero.wall_tracer.trackDistX[-8] ),
    .A1(_09844_),
    .S(_05414_),
    .X(_09845_));
 sky130_fd_sc_hd__clkbuf_1 _17271_ (.A(_09845_),
    .X(_00581_));
 sky130_fd_sc_hd__or2_1 _17272_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .X(_09846_));
 sky130_fd_sc_hd__nand2_1 _17273_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09847_));
 sky130_fd_sc_hd__o21bai_2 _17274_ (.A1(_09838_),
    .A2(_09840_),
    .B1_N(_09839_),
    .Y(_09848_));
 sky130_fd_sc_hd__and3_1 _17275_ (.A(_09846_),
    .B(_09847_),
    .C(_09848_),
    .X(_09849_));
 sky130_fd_sc_hd__a21oi_1 _17276_ (.A1(_09846_),
    .A2(_09847_),
    .B1(_09848_),
    .Y(_09850_));
 sky130_fd_sc_hd__nand2_1 _17277_ (.A(_05531_),
    .B(_09076_),
    .Y(_09851_));
 sky130_fd_sc_hd__o31ai_1 _17278_ (.A1(_09812_),
    .A2(_09849_),
    .A3(_09850_),
    .B1(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__mux2_1 _17279_ (.A0(\rbzero.wall_tracer.trackDistX[-7] ),
    .A1(_09852_),
    .S(_05413_),
    .X(_09853_));
 sky130_fd_sc_hd__clkbuf_1 _17280_ (.A(_09853_),
    .X(_00582_));
 sky130_fd_sc_hd__nor2_1 _17281_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_09854_));
 sky130_fd_sc_hd__and2_1 _17282_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_09855_));
 sky130_fd_sc_hd__a21boi_1 _17283_ (.A1(_09846_),
    .A2(_09848_),
    .B1_N(_09847_),
    .Y(_09856_));
 sky130_fd_sc_hd__nor3_1 _17284_ (.A(_09854_),
    .B(_09855_),
    .C(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__o21a_1 _17285_ (.A1(_09854_),
    .A2(_09855_),
    .B1(_09856_),
    .X(_09858_));
 sky130_fd_sc_hd__nand2_2 _17286_ (.A(_09061_),
    .B(_09062_),
    .Y(_09859_));
 sky130_fd_sc_hd__or2_1 _17287_ (.A(_09807_),
    .B(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__o31ai_1 _17288_ (.A1(_09812_),
    .A2(_09857_),
    .A3(_09858_),
    .B1(_09860_),
    .Y(_09861_));
 sky130_fd_sc_hd__mux2_1 _17289_ (.A0(\rbzero.wall_tracer.trackDistX[-6] ),
    .A1(_09861_),
    .S(_05413_),
    .X(_09862_));
 sky130_fd_sc_hd__clkbuf_1 _17290_ (.A(_09862_),
    .X(_00583_));
 sky130_fd_sc_hd__buf_4 _17291_ (.A(_04016_),
    .X(_09863_));
 sky130_fd_sc_hd__or2_1 _17292_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .X(_09864_));
 sky130_fd_sc_hd__nand2_1 _17293_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09865_));
 sky130_fd_sc_hd__o21bai_1 _17294_ (.A1(_09854_),
    .A2(_09856_),
    .B1_N(_09855_),
    .Y(_09866_));
 sky130_fd_sc_hd__and3_1 _17295_ (.A(_09864_),
    .B(_09865_),
    .C(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__a21oi_1 _17296_ (.A1(_09864_),
    .A2(_09865_),
    .B1(_09866_),
    .Y(_09868_));
 sky130_fd_sc_hd__or2_1 _17297_ (.A(_09807_),
    .B(_09194_),
    .X(_09869_));
 sky130_fd_sc_hd__o31ai_1 _17298_ (.A1(_09863_),
    .A2(_09867_),
    .A3(_09868_),
    .B1(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__mux2_1 _17299_ (.A0(\rbzero.wall_tracer.trackDistX[-5] ),
    .A1(_09870_),
    .S(_05413_),
    .X(_09871_));
 sky130_fd_sc_hd__clkbuf_1 _17300_ (.A(_09871_),
    .X(_00584_));
 sky130_fd_sc_hd__nor2_1 _17301_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09872_));
 sky130_fd_sc_hd__nand2_1 _17302_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09873_));
 sky130_fd_sc_hd__or2b_1 _17303_ (.A(_09872_),
    .B_N(_09873_),
    .X(_09874_));
 sky130_fd_sc_hd__a21boi_1 _17304_ (.A1(_09864_),
    .A2(_09866_),
    .B1_N(_09865_),
    .Y(_09875_));
 sky130_fd_sc_hd__xnor2_1 _17305_ (.A(_09874_),
    .B(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__or2_1 _17306_ (.A(_09807_),
    .B(_09331_),
    .X(_09877_));
 sky130_fd_sc_hd__o21ai_1 _17307_ (.A1(_09812_),
    .A2(_09876_),
    .B1(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__mux2_1 _17308_ (.A0(\rbzero.wall_tracer.trackDistX[-4] ),
    .A1(_09878_),
    .S(_05413_),
    .X(_09879_));
 sky130_fd_sc_hd__clkbuf_1 _17309_ (.A(_09879_),
    .X(_00585_));
 sky130_fd_sc_hd__or2_1 _17310_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .X(_09880_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09881_));
 sky130_fd_sc_hd__o21ai_1 _17312_ (.A1(_09872_),
    .A2(_09875_),
    .B1(_09873_),
    .Y(_09882_));
 sky130_fd_sc_hd__and3_1 _17313_ (.A(_09880_),
    .B(_09881_),
    .C(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__a21oi_1 _17314_ (.A1(_09880_),
    .A2(_09881_),
    .B1(_09882_),
    .Y(_09884_));
 sky130_fd_sc_hd__or2_1 _17315_ (.A(_09807_),
    .B(_09458_),
    .X(_09885_));
 sky130_fd_sc_hd__o31ai_1 _17316_ (.A1(_09863_),
    .A2(_09883_),
    .A3(_09884_),
    .B1(_09885_),
    .Y(_09886_));
 sky130_fd_sc_hd__mux2_1 _17317_ (.A0(\rbzero.wall_tracer.trackDistX[-3] ),
    .A1(_09886_),
    .S(_05413_),
    .X(_09887_));
 sky130_fd_sc_hd__clkbuf_1 _17318_ (.A(_09887_),
    .X(_00586_));
 sky130_fd_sc_hd__and2_1 _17319_ (.A(_05532_),
    .B(_09597_),
    .X(_09888_));
 sky130_fd_sc_hd__clkbuf_4 _17320_ (.A(_05394_),
    .X(_09889_));
 sky130_fd_sc_hd__nor2_1 _17321_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09890_));
 sky130_fd_sc_hd__and2_1 _17322_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_09891_));
 sky130_fd_sc_hd__a21boi_1 _17323_ (.A1(_09880_),
    .A2(_09882_),
    .B1_N(_09881_),
    .Y(_09892_));
 sky130_fd_sc_hd__or3_1 _17324_ (.A(_09890_),
    .B(_09891_),
    .C(_09892_),
    .X(_09893_));
 sky130_fd_sc_hd__o21ai_1 _17325_ (.A1(_09890_),
    .A2(_09891_),
    .B1(_09892_),
    .Y(_09894_));
 sky130_fd_sc_hd__a31o_1 _17326_ (.A1(_09889_),
    .A2(_09893_),
    .A3(_09894_),
    .B1(_09780_),
    .X(_09895_));
 sky130_fd_sc_hd__o22a_1 _17327_ (.A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .A2(_09817_),
    .B1(_09888_),
    .B2(_09895_),
    .X(_00587_));
 sky130_fd_sc_hd__nand2_1 _17328_ (.A(_04016_),
    .B(_09739_),
    .Y(_09896_));
 sky130_fd_sc_hd__inv_2 _17329_ (.A(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__nor2_1 _17330_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_09898_));
 sky130_fd_sc_hd__and2_1 _17331_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_09899_));
 sky130_fd_sc_hd__nand2_1 _17332_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09900_));
 sky130_fd_sc_hd__o211ai_1 _17333_ (.A1(_09898_),
    .A2(_09899_),
    .B1(_09900_),
    .C1(_09893_),
    .Y(_09901_));
 sky130_fd_sc_hd__a211o_1 _17334_ (.A1(_09900_),
    .A2(_09893_),
    .B1(_09898_),
    .C1(_09899_),
    .X(_09902_));
 sky130_fd_sc_hd__a31o_1 _17335_ (.A1(_09889_),
    .A2(_09901_),
    .A3(_09902_),
    .B1(_09780_),
    .X(_09903_));
 sky130_fd_sc_hd__o22a_1 _17336_ (.A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .A2(_09817_),
    .B1(_09897_),
    .B2(_09903_),
    .X(_00588_));
 sky130_fd_sc_hd__or3_1 _17337_ (.A(_09605_),
    .B(_09606_),
    .C(_09734_),
    .X(_09904_));
 sky130_fd_sc_hd__a21o_1 _17338_ (.A1(_09592_),
    .A2(_09904_),
    .B1(_09736_),
    .X(_09905_));
 sky130_fd_sc_hd__a31oi_4 _17339_ (.A1(_09594_),
    .A2(_09596_),
    .A3(_09737_),
    .B1(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__and2b_1 _17340_ (.A_N(_09486_),
    .B(_09495_),
    .X(_09907_));
 sky130_fd_sc_hd__a21o_2 _17341_ (.A1(_09609_),
    .A2(_09612_),
    .B1(_09907_),
    .X(_09908_));
 sky130_fd_sc_hd__or2b_1 _17342_ (.A(_09656_),
    .B_N(_09617_),
    .X(_09909_));
 sky130_fd_sc_hd__nand2_1 _17343_ (.A(_08331_),
    .B(_09621_),
    .Y(_09910_));
 sky130_fd_sc_hd__o31a_1 _17344_ (.A1(_08335_),
    .A2(_09359_),
    .A3(_09910_),
    .B1(_09624_),
    .X(_09911_));
 sky130_fd_sc_hd__a21oi_2 _17345_ (.A1(_09633_),
    .A2(_09636_),
    .B1(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__and3_1 _17346_ (.A(_09633_),
    .B(_09636_),
    .C(_09911_),
    .X(_09913_));
 sky130_fd_sc_hd__or2_1 _17347_ (.A(_09912_),
    .B(_09913_),
    .X(_09914_));
 sky130_fd_sc_hd__a21oi_1 _17348_ (.A1(_09654_),
    .A2(_09909_),
    .B1(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__and3_1 _17349_ (.A(_09654_),
    .B(_09909_),
    .C(_09914_),
    .X(_09916_));
 sky130_fd_sc_hd__nor2_2 _17350_ (.A(_09915_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__xor2_4 _17351_ (.A(_09908_),
    .B(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__a21o_1 _17352_ (.A1(_09638_),
    .A2(_09652_),
    .B1(_09650_),
    .X(_09919_));
 sky130_fd_sc_hd__or2b_1 _17353_ (.A(_09678_),
    .B_N(_09660_),
    .X(_09920_));
 sky130_fd_sc_hd__or2b_1 _17354_ (.A(_09679_),
    .B_N(_09659_),
    .X(_09921_));
 sky130_fd_sc_hd__or3_1 _17355_ (.A(_08335_),
    .B(_09483_),
    .C(_09910_),
    .X(_09922_));
 sky130_fd_sc_hd__o21ai_1 _17356_ (.A1(_08335_),
    .A2(_09483_),
    .B1(_09910_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_1 _17357_ (.A(_09922_),
    .B(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__nor2_1 _17358_ (.A(_08416_),
    .B(_09704_),
    .Y(_09925_));
 sky130_fd_sc_hd__xnor2_1 _17359_ (.A(_09924_),
    .B(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__or4_1 _17360_ (.A(_09243_),
    .B(_08821_),
    .C(_09028_),
    .D(_09164_),
    .X(_09927_));
 sky130_fd_sc_hd__o22ai_1 _17361_ (.A1(_09243_),
    .A2(_09029_),
    .B1(_09164_),
    .B2(_09096_),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_1 _17362_ (.A(_09927_),
    .B(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__nor2_1 _17363_ (.A(_09368_),
    .B(_09217_),
    .Y(_09930_));
 sky130_fd_sc_hd__xor2_1 _17364_ (.A(_09929_),
    .B(_09930_),
    .X(_09931_));
 sky130_fd_sc_hd__o31a_1 _17365_ (.A1(_09368_),
    .A2(_09165_),
    .A3(_09628_),
    .B1(_09629_),
    .X(_09932_));
 sky130_fd_sc_hd__or2_1 _17366_ (.A(_09931_),
    .B(_09932_),
    .X(_09933_));
 sky130_fd_sc_hd__nand2_1 _17367_ (.A(_09931_),
    .B(_09932_),
    .Y(_09934_));
 sky130_fd_sc_hd__and2_1 _17368_ (.A(_09933_),
    .B(_09934_),
    .X(_09935_));
 sky130_fd_sc_hd__nand2_1 _17369_ (.A(_09926_),
    .B(_09935_),
    .Y(_09936_));
 sky130_fd_sc_hd__or2_1 _17370_ (.A(_09926_),
    .B(_09935_),
    .X(_09937_));
 sky130_fd_sc_hd__and2_1 _17371_ (.A(_09936_),
    .B(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__a21bo_1 _17372_ (.A1(_09641_),
    .A2(_09644_),
    .B1_N(_09643_),
    .X(_09939_));
 sky130_fd_sc_hd__nand2_1 _17373_ (.A(_09664_),
    .B(_09665_),
    .Y(_09940_));
 sky130_fd_sc_hd__o22a_1 _17374_ (.A1(_08705_),
    .A2(_08159_),
    .B1(_08151_),
    .B2(_09522_),
    .X(_09941_));
 sky130_fd_sc_hd__or3_1 _17375_ (.A(_09522_),
    .B(_08705_),
    .C(_08419_),
    .X(_09942_));
 sky130_fd_sc_hd__or2b_1 _17376_ (.A(_09941_),
    .B_N(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__nor2_1 _17377_ (.A(_09245_),
    .B(_08427_),
    .Y(_09944_));
 sky130_fd_sc_hd__xor2_1 _17378_ (.A(_09943_),
    .B(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__xnor2_1 _17379_ (.A(_09940_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__xnor2_1 _17380_ (.A(_09939_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__a21oi_1 _17381_ (.A1(_09521_),
    .A2(_09525_),
    .B1(_09645_),
    .Y(_09948_));
 sky130_fd_sc_hd__a21oi_2 _17382_ (.A1(_09639_),
    .A2(_09646_),
    .B1(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__xor2_1 _17383_ (.A(_09947_),
    .B(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__xnor2_1 _17384_ (.A(_09938_),
    .B(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__a21o_1 _17385_ (.A1(_09920_),
    .A2(_09921_),
    .B1(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__nand3_1 _17386_ (.A(_09920_),
    .B(_09921_),
    .C(_09951_),
    .Y(_09953_));
 sky130_fd_sc_hd__nand2_1 _17387_ (.A(_09952_),
    .B(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__xnor2_2 _17388_ (.A(_09919_),
    .B(_09954_),
    .Y(_09955_));
 sky130_fd_sc_hd__nor2_1 _17389_ (.A(_09673_),
    .B(_09676_),
    .Y(_09956_));
 sky130_fd_sc_hd__a31o_1 _17390_ (.A1(_09665_),
    .A2(_09666_),
    .A3(_09677_),
    .B1(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__a21o_2 _17391_ (.A1(_09682_),
    .A2(_09690_),
    .B1(_09689_),
    .X(_09958_));
 sky130_fd_sc_hd__nand2_1 _17392_ (.A(_08445_),
    .B(_08332_),
    .Y(_09959_));
 sky130_fd_sc_hd__xnor2_1 _17393_ (.A(_09663_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__or3_1 _17394_ (.A(_09661_),
    .B(_08356_),
    .C(_09960_),
    .X(_09961_));
 sky130_fd_sc_hd__o21ai_1 _17395_ (.A1(_09661_),
    .A2(_08356_),
    .B1(_09960_),
    .Y(_09962_));
 sky130_fd_sc_hd__and2_1 _17396_ (.A(_09961_),
    .B(_09962_),
    .X(_09963_));
 sky130_fd_sc_hd__nor2_1 _17397_ (.A(_09126_),
    .B(_08570_),
    .Y(_09964_));
 sky130_fd_sc_hd__xnor2_2 _17398_ (.A(_09670_),
    .B(_09964_),
    .Y(_09965_));
 sky130_fd_sc_hd__or2_1 _17399_ (.A(_08178_),
    .B(_09103_),
    .X(_09966_));
 sky130_fd_sc_hd__xnor2_2 _17400_ (.A(_09965_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__a22oi_4 _17401_ (.A1(_09545_),
    .A2(_09670_),
    .B1(_09672_),
    .B2(_09669_),
    .Y(_09968_));
 sky130_fd_sc_hd__xor2_2 _17402_ (.A(_09967_),
    .B(_09968_),
    .X(_09969_));
 sky130_fd_sc_hd__xor2_2 _17403_ (.A(_09963_),
    .B(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__xnor2_1 _17404_ (.A(_09958_),
    .B(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__xnor2_1 _17405_ (.A(_09957_),
    .B(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__clkbuf_4 _17406_ (.A(_09540_),
    .X(_09973_));
 sky130_fd_sc_hd__nor2_1 _17407_ (.A(_08895_),
    .B(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__a22o_1 _17408_ (.A1(_09553_),
    .A2(_09974_),
    .B1(_09687_),
    .B2(_09684_),
    .X(_09975_));
 sky130_fd_sc_hd__and2_1 _17409_ (.A(_09288_),
    .B(_09695_),
    .X(_09976_));
 sky130_fd_sc_hd__clkbuf_4 _17410_ (.A(_09976_),
    .X(_09977_));
 sky130_fd_sc_hd__or3_1 _17411_ (.A(_08872_),
    .B(_09977_),
    .C(_09700_),
    .X(_09978_));
 sky130_fd_sc_hd__a21bo_1 _17412_ (.A1(_09694_),
    .A2(_09701_),
    .B1_N(_09978_),
    .X(_09979_));
 sky130_fd_sc_hd__nor2_2 _17413_ (.A(_08284_),
    .B(_09540_),
    .Y(_09980_));
 sky130_fd_sc_hd__o22a_1 _17414_ (.A1(_08767_),
    .A2(_09552_),
    .B1(_09973_),
    .B2(_08283_),
    .X(_09981_));
 sky130_fd_sc_hd__a21o_1 _17415_ (.A1(_09686_),
    .A2(_09980_),
    .B1(_09981_),
    .X(_09982_));
 sky130_fd_sc_hd__nor2_1 _17416_ (.A(_09114_),
    .B(_09417_),
    .Y(_09983_));
 sky130_fd_sc_hd__xnor2_2 _17417_ (.A(_09982_),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__xor2_2 _17418_ (.A(_09979_),
    .B(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__xor2_2 _17419_ (.A(_09975_),
    .B(_09985_),
    .X(_09986_));
 sky130_fd_sc_hd__nor2_1 _17420_ (.A(_09117_),
    .B(_09693_),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_1 _17421_ (.A(_05210_),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_09988_));
 sky130_fd_sc_hd__nand2_1 _17422_ (.A(_09434_),
    .B(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__and2_1 _17423_ (.A(_09434_),
    .B(_09988_),
    .X(_09990_));
 sky130_fd_sc_hd__clkbuf_4 _17424_ (.A(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__o22a_1 _17425_ (.A1(_08873_),
    .A2(_09977_),
    .B1(_09991_),
    .B2(_08872_),
    .X(_09992_));
 sky130_fd_sc_hd__a31oi_2 _17426_ (.A1(_08266_),
    .A2(_09696_),
    .A3(_09989_),
    .B1(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__xor2_2 _17427_ (.A(_09987_),
    .B(_09993_),
    .X(_09994_));
 sky130_fd_sc_hd__or3_1 _17428_ (.A(_05211_),
    .B(_08215_),
    .C(_09565_),
    .X(_09995_));
 sky130_fd_sc_hd__or2_1 _17429_ (.A(_08519_),
    .B(_09699_),
    .X(_09996_));
 sky130_fd_sc_hd__mux2_1 _17430_ (.A0(_07601_),
    .A1(_09995_),
    .S(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__a21o_1 _17431_ (.A1(_08377_),
    .A2(_08519_),
    .B1(_09699_),
    .X(_09998_));
 sky130_fd_sc_hd__o21ai_1 _17432_ (.A1(_08747_),
    .A2(_09699_),
    .B1(_08250_),
    .Y(_09999_));
 sky130_fd_sc_hd__o2bb2a_2 _17433_ (.A1_N(_09700_),
    .A2_N(_09997_),
    .B1(_09998_),
    .B2(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__o21a_1 _17434_ (.A1(_09707_),
    .A2(_09708_),
    .B1(_09706_),
    .X(_10001_));
 sky130_fd_sc_hd__xnor2_2 _17435_ (.A(_10000_),
    .B(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__xnor2_1 _17436_ (.A(_09994_),
    .B(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__nor2_1 _17437_ (.A(_09709_),
    .B(_09712_),
    .Y(_10004_));
 sky130_fd_sc_hd__a21o_1 _17438_ (.A1(_09702_),
    .A2(_09713_),
    .B1(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__xnor2_2 _17439_ (.A(_10003_),
    .B(_10005_),
    .Y(_10006_));
 sky130_fd_sc_hd__xnor2_2 _17440_ (.A(_09986_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__nor2_1 _17441_ (.A(_09714_),
    .B(_09716_),
    .Y(_10008_));
 sky130_fd_sc_hd__a21o_2 _17442_ (.A1(_09692_),
    .A2(_09717_),
    .B1(_10008_),
    .X(_10009_));
 sky130_fd_sc_hd__xnor2_1 _17443_ (.A(_10007_),
    .B(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__xnor2_1 _17444_ (.A(_09972_),
    .B(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__nor2_1 _17445_ (.A(_09718_),
    .B(_09720_),
    .Y(_10012_));
 sky130_fd_sc_hd__a21o_1 _17446_ (.A1(_09680_),
    .A2(_09721_),
    .B1(_10012_),
    .X(_10013_));
 sky130_fd_sc_hd__xnor2_1 _17447_ (.A(_10011_),
    .B(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__xnor2_2 _17448_ (.A(_09955_),
    .B(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__nor2_1 _17449_ (.A(_09722_),
    .B(_09724_),
    .Y(_10016_));
 sky130_fd_sc_hd__a21o_1 _17450_ (.A1(_09657_),
    .A2(_09725_),
    .B1(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__xnor2_2 _17451_ (.A(_10015_),
    .B(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__xnor2_4 _17452_ (.A(_09918_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__nor2_1 _17453_ (.A(_09726_),
    .B(_09728_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21oi_2 _17454_ (.A1(_09616_),
    .A2(_09729_),
    .B1(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__xor2_4 _17455_ (.A(_10019_),
    .B(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__xnor2_4 _17456_ (.A(_09614_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__nor2_1 _17457_ (.A(_09730_),
    .B(_09732_),
    .Y(_10024_));
 sky130_fd_sc_hd__a21oi_4 _17458_ (.A1(_09474_),
    .A2(_09733_),
    .B1(_10024_),
    .Y(_10025_));
 sky130_fd_sc_hd__xor2_4 _17459_ (.A(_10023_),
    .B(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__xor2_4 _17460_ (.A(_09906_),
    .B(_10026_),
    .X(_10027_));
 sky130_fd_sc_hd__or2_1 _17461_ (.A(_09889_),
    .B(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__nand2_1 _17462_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_10029_));
 sky130_fd_sc_hd__nor2_1 _17463_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_10030_));
 sky130_fd_sc_hd__and2_1 _17464_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_10031_));
 sky130_fd_sc_hd__a211o_1 _17465_ (.A1(_10029_),
    .A2(_09902_),
    .B1(_10030_),
    .C1(_10031_),
    .X(_10032_));
 sky130_fd_sc_hd__inv_2 _17466_ (.A(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__o211a_1 _17467_ (.A1(_10030_),
    .A2(_10031_),
    .B1(_10029_),
    .C1(_09902_),
    .X(_10034_));
 sky130_fd_sc_hd__o31a_1 _17468_ (.A1(_05532_),
    .A2(_10033_),
    .A3(_10034_),
    .B1(_09817_),
    .X(_10035_));
 sky130_fd_sc_hd__buf_2 _17469_ (.A(_09817_),
    .X(_10036_));
 sky130_fd_sc_hd__o2bb2a_1 _17470_ (.A1_N(_10028_),
    .A2_N(_10035_),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_10036_),
    .X(_00589_));
 sky130_fd_sc_hd__or2_1 _17471_ (.A(_10019_),
    .B(_10021_),
    .X(_10037_));
 sky130_fd_sc_hd__nand2_1 _17472_ (.A(_09614_),
    .B(_10022_),
    .Y(_10038_));
 sky130_fd_sc_hd__a21o_1 _17473_ (.A1(_09908_),
    .A2(_09917_),
    .B1(_09915_),
    .X(_10039_));
 sky130_fd_sc_hd__or2b_1 _17474_ (.A(_09954_),
    .B_N(_09919_),
    .X(_10040_));
 sky130_fd_sc_hd__o31a_1 _17475_ (.A1(_08416_),
    .A2(_09704_),
    .A3(_09924_),
    .B1(_09922_),
    .X(_10041_));
 sky130_fd_sc_hd__a21oi_2 _17476_ (.A1(_09933_),
    .A2(_09936_),
    .B1(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__and3_1 _17477_ (.A(_09933_),
    .B(_09936_),
    .C(_10041_),
    .X(_10043_));
 sky130_fd_sc_hd__or2_1 _17478_ (.A(_10042_),
    .B(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__a21oi_1 _17479_ (.A1(_09952_),
    .A2(_10040_),
    .B1(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__and3_1 _17480_ (.A(_09952_),
    .B(_10040_),
    .C(_10044_),
    .X(_10046_));
 sky130_fd_sc_hd__nor2_1 _17481_ (.A(_10045_),
    .B(_10046_),
    .Y(_10047_));
 sky130_fd_sc_hd__xor2_1 _17482_ (.A(_09912_),
    .B(_10047_),
    .X(_10048_));
 sky130_fd_sc_hd__nor2_1 _17483_ (.A(_09947_),
    .B(_09949_),
    .Y(_10049_));
 sky130_fd_sc_hd__a21o_1 _17484_ (.A1(_09938_),
    .A2(_09950_),
    .B1(_10049_),
    .X(_10050_));
 sky130_fd_sc_hd__nand2_1 _17485_ (.A(_09958_),
    .B(_09970_),
    .Y(_10051_));
 sky130_fd_sc_hd__or2b_1 _17486_ (.A(_09971_),
    .B_N(_09957_),
    .X(_10052_));
 sky130_fd_sc_hd__o22ai_1 _17487_ (.A1(_09368_),
    .A2(_09480_),
    .B1(_09483_),
    .B2(_08329_),
    .Y(_10053_));
 sky130_fd_sc_hd__or3_1 _17488_ (.A(_09368_),
    .B(_09483_),
    .C(_09910_),
    .X(_10054_));
 sky130_fd_sc_hd__nand2_1 _17489_ (.A(_10053_),
    .B(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__and2_1 _17490_ (.A(_08335_),
    .B(_09703_),
    .X(_10056_));
 sky130_fd_sc_hd__xnor2_1 _17491_ (.A(_10055_),
    .B(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__o22ai_1 _17492_ (.A1(_09245_),
    .A2(_09029_),
    .B1(_09165_),
    .B2(_09243_),
    .Y(_10058_));
 sky130_fd_sc_hd__or4_1 _17493_ (.A(_09245_),
    .B(_09243_),
    .C(_09028_),
    .D(_09164_),
    .X(_10059_));
 sky130_fd_sc_hd__nand2_1 _17494_ (.A(_10058_),
    .B(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__nor2_1 _17495_ (.A(_09096_),
    .B(_09217_),
    .Y(_10061_));
 sky130_fd_sc_hd__xor2_1 _17496_ (.A(_10060_),
    .B(_10061_),
    .X(_10062_));
 sky130_fd_sc_hd__o31a_1 _17497_ (.A1(_09368_),
    .A2(_09217_),
    .A3(_09929_),
    .B1(_09927_),
    .X(_10063_));
 sky130_fd_sc_hd__or2_1 _17498_ (.A(_10062_),
    .B(_10063_),
    .X(_10064_));
 sky130_fd_sc_hd__nand2_1 _17499_ (.A(_10062_),
    .B(_10063_),
    .Y(_10065_));
 sky130_fd_sc_hd__and2_1 _17500_ (.A(_10064_),
    .B(_10065_),
    .X(_10066_));
 sky130_fd_sc_hd__nand2_1 _17501_ (.A(_10057_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__or2_1 _17502_ (.A(_10057_),
    .B(_10066_),
    .X(_10068_));
 sky130_fd_sc_hd__and2_1 _17503_ (.A(_10067_),
    .B(_10068_),
    .X(_10069_));
 sky130_fd_sc_hd__o31ai_2 _17504_ (.A1(_09391_),
    .A2(_08427_),
    .A3(_09941_),
    .B1(_09942_),
    .Y(_10070_));
 sky130_fd_sc_hd__or2_1 _17505_ (.A(_09663_),
    .B(_09959_),
    .X(_10071_));
 sky130_fd_sc_hd__nand2_1 _17506_ (.A(_10071_),
    .B(_09961_),
    .Y(_10072_));
 sky130_fd_sc_hd__o22ai_1 _17507_ (.A1(_09522_),
    .A2(_08159_),
    .B1(_08151_),
    .B2(_09661_),
    .Y(_10073_));
 sky130_fd_sc_hd__or2_1 _17508_ (.A(_07974_),
    .B(_08158_),
    .X(_10074_));
 sky130_fd_sc_hd__or3_1 _17509_ (.A(_09522_),
    .B(_08151_),
    .C(_10074_),
    .X(_10075_));
 sky130_fd_sc_hd__nand2_1 _17510_ (.A(_10073_),
    .B(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__nor2_1 _17511_ (.A(_09526_),
    .B(_08427_),
    .Y(_10077_));
 sky130_fd_sc_hd__xor2_1 _17512_ (.A(_10076_),
    .B(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__xnor2_1 _17513_ (.A(_10072_),
    .B(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__xnor2_1 _17514_ (.A(_10070_),
    .B(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__a21oi_1 _17515_ (.A1(_09664_),
    .A2(_09665_),
    .B1(_09945_),
    .Y(_10081_));
 sky130_fd_sc_hd__a21oi_1 _17516_ (.A1(_09939_),
    .A2(_09946_),
    .B1(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__xor2_1 _17517_ (.A(_10080_),
    .B(_10082_),
    .X(_10083_));
 sky130_fd_sc_hd__xnor2_1 _17518_ (.A(_10069_),
    .B(_10083_),
    .Y(_10084_));
 sky130_fd_sc_hd__a21o_1 _17519_ (.A1(_10051_),
    .A2(_10052_),
    .B1(_10084_),
    .X(_10085_));
 sky130_fd_sc_hd__nand3_1 _17520_ (.A(_10051_),
    .B(_10052_),
    .C(_10084_),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_1 _17521_ (.A(_10085_),
    .B(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__xnor2_1 _17522_ (.A(_10050_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__nor2_1 _17523_ (.A(_09967_),
    .B(_09968_),
    .Y(_10089_));
 sky130_fd_sc_hd__a21o_1 _17524_ (.A1(_09963_),
    .A2(_09969_),
    .B1(_10089_),
    .X(_10090_));
 sky130_fd_sc_hd__and2_1 _17525_ (.A(_09979_),
    .B(_09984_),
    .X(_10091_));
 sky130_fd_sc_hd__a21oi_2 _17526_ (.A1(_09975_),
    .A2(_09985_),
    .B1(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__or4_1 _17527_ (.A(_08178_),
    .B(_08202_),
    .C(_08493_),
    .D(_08044_),
    .X(_10093_));
 sky130_fd_sc_hd__clkbuf_4 _17528_ (.A(_08202_),
    .X(_10094_));
 sky130_fd_sc_hd__o22ai_1 _17529_ (.A1(_08178_),
    .A2(_08493_),
    .B1(_08044_),
    .B2(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__nand2_1 _17530_ (.A(_10093_),
    .B(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__nor2_1 _17531_ (.A(_08275_),
    .B(_08356_),
    .Y(_10097_));
 sky130_fd_sc_hd__xnor2_2 _17532_ (.A(_10096_),
    .B(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__nor2_2 _17533_ (.A(_09668_),
    .B(_09417_),
    .Y(_10099_));
 sky130_fd_sc_hd__o22a_1 _17534_ (.A1(_09276_),
    .A2(_08570_),
    .B1(_09417_),
    .B2(_08111_),
    .X(_10100_));
 sky130_fd_sc_hd__a21o_1 _17535_ (.A1(_09670_),
    .A2(_10099_),
    .B1(_10100_),
    .X(_10101_));
 sky130_fd_sc_hd__nor2_1 _17536_ (.A(_09126_),
    .B(_09674_),
    .Y(_10102_));
 sky130_fd_sc_hd__xor2_2 _17537_ (.A(_10101_),
    .B(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__nand2_1 _17538_ (.A(_09670_),
    .B(_09964_),
    .Y(_10104_));
 sky130_fd_sc_hd__o31a_1 _17539_ (.A1(_08178_),
    .A2(_09674_),
    .A3(_09965_),
    .B1(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__xor2_2 _17540_ (.A(_10103_),
    .B(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__xnor2_2 _17541_ (.A(_10098_),
    .B(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__xor2_2 _17542_ (.A(_10092_),
    .B(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__xor2_2 _17543_ (.A(_10090_),
    .B(_10108_),
    .X(_10109_));
 sky130_fd_sc_hd__clkbuf_4 _17544_ (.A(_09114_),
    .X(_10110_));
 sky130_fd_sc_hd__or3_1 _17545_ (.A(_10110_),
    .B(_09417_),
    .C(_09982_),
    .X(_10111_));
 sky130_fd_sc_hd__a21bo_1 _17546_ (.A1(_09686_),
    .A2(_09980_),
    .B1_N(_10111_),
    .X(_10112_));
 sky130_fd_sc_hd__or3b_1 _17547_ (.A(_08873_),
    .B(_09991_),
    .C_N(_09696_),
    .X(_10113_));
 sky130_fd_sc_hd__o31a_1 _17548_ (.A1(_09117_),
    .A2(_09693_),
    .A3(_09992_),
    .B1(_10113_),
    .X(_10114_));
 sky130_fd_sc_hd__nor2_1 _17549_ (.A(_08283_),
    .B(_09555_),
    .Y(_10115_));
 sky130_fd_sc_hd__xnor2_1 _17550_ (.A(_09980_),
    .B(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__nor2_1 _17551_ (.A(_09114_),
    .B(_09552_),
    .Y(_10117_));
 sky130_fd_sc_hd__xnor2_1 _17552_ (.A(_10116_),
    .B(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__and2b_1 _17553_ (.A_N(_10114_),
    .B(_10118_),
    .X(_10119_));
 sky130_fd_sc_hd__or2b_1 _17554_ (.A(_10118_),
    .B_N(_10114_),
    .X(_10120_));
 sky130_fd_sc_hd__or2b_1 _17555_ (.A(_10119_),
    .B_N(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__xnor2_2 _17556_ (.A(_10112_),
    .B(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__or2b_1 _17557_ (.A(_10001_),
    .B_N(_10000_),
    .X(_10123_));
 sky130_fd_sc_hd__a21bo_1 _17558_ (.A1(_09994_),
    .A2(_10002_),
    .B1_N(_10123_),
    .X(_10124_));
 sky130_fd_sc_hd__nor2_1 _17559_ (.A(_08747_),
    .B(_09700_),
    .Y(_10125_));
 sky130_fd_sc_hd__and2_1 _17560_ (.A(_09700_),
    .B(_09998_),
    .X(_10126_));
 sky130_fd_sc_hd__or2_1 _17561_ (.A(_10125_),
    .B(_10126_),
    .X(_10127_));
 sky130_fd_sc_hd__nand2_2 _17562_ (.A(_05211_),
    .B(\rbzero.wall_tracer.stepDistX[11] ),
    .Y(_10128_));
 sky130_fd_sc_hd__o21a_1 _17563_ (.A1(_05211_),
    .A2(_09699_),
    .B1(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__or3_1 _17564_ (.A(_08872_),
    .B(_08873_),
    .C(_10129_),
    .X(_10130_));
 sky130_fd_sc_hd__nand2_1 _17565_ (.A(_08872_),
    .B(_08873_),
    .Y(_10131_));
 sky130_fd_sc_hd__nor2_1 _17566_ (.A(_09117_),
    .B(_10129_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand3_1 _17567_ (.A(_10130_),
    .B(_10131_),
    .C(_10132_),
    .Y(_10133_));
 sky130_fd_sc_hd__o21ai_2 _17568_ (.A1(_05211_),
    .A2(_09699_),
    .B1(_10128_),
    .Y(_10134_));
 sky130_fd_sc_hd__a31o_1 _17569_ (.A1(_10134_),
    .A2(_10130_),
    .A3(_10131_),
    .B1(_10132_),
    .X(_10135_));
 sky130_fd_sc_hd__and2_1 _17570_ (.A(_10133_),
    .B(_10135_),
    .X(_10136_));
 sky130_fd_sc_hd__nor2_1 _17571_ (.A(_09117_),
    .B(_09977_),
    .Y(_10137_));
 sky130_fd_sc_hd__inv_2 _17572_ (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_10138_));
 sky130_fd_sc_hd__mux2_4 _17573_ (.A0(_10138_),
    .A1(_09565_),
    .S(_05198_),
    .X(_10139_));
 sky130_fd_sc_hd__or4_1 _17574_ (.A(_08872_),
    .B(_08873_),
    .C(_09991_),
    .D(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__a2bb2o_1 _17575_ (.A1_N(_08872_),
    .A2_N(_10139_),
    .B1(_08266_),
    .B2(_09989_),
    .X(_10141_));
 sky130_fd_sc_hd__and3_1 _17576_ (.A(_10137_),
    .B(_10140_),
    .C(_10141_),
    .X(_10142_));
 sky130_fd_sc_hd__a21o_1 _17577_ (.A1(_10140_),
    .A2(_10141_),
    .B1(_10137_),
    .X(_10143_));
 sky130_fd_sc_hd__nand2_1 _17578_ (.A(_10127_),
    .B(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__o22a_1 _17579_ (.A1(_10127_),
    .A2(_10136_),
    .B1(_10142_),
    .B2(_10144_),
    .X(_10145_));
 sky130_fd_sc_hd__xnor2_2 _17580_ (.A(_10124_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__xnor2_2 _17581_ (.A(_10122_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__nand2_1 _17582_ (.A(_09994_),
    .B(_10002_),
    .Y(_10148_));
 sky130_fd_sc_hd__or2_1 _17583_ (.A(_09994_),
    .B(_10002_),
    .X(_10149_));
 sky130_fd_sc_hd__a32o_2 _17584_ (.A1(_10148_),
    .A2(_10149_),
    .A3(_10005_),
    .B1(_10006_),
    .B2(_09986_),
    .X(_10150_));
 sky130_fd_sc_hd__xnor2_1 _17585_ (.A(_10147_),
    .B(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__xnor2_1 _17586_ (.A(_10109_),
    .B(_10151_),
    .Y(_10152_));
 sky130_fd_sc_hd__or2b_1 _17587_ (.A(_10007_),
    .B_N(_10009_),
    .X(_10153_));
 sky130_fd_sc_hd__a21boi_1 _17588_ (.A1(_09972_),
    .A2(_10010_),
    .B1_N(_10153_),
    .Y(_10154_));
 sky130_fd_sc_hd__xor2_1 _17589_ (.A(_10152_),
    .B(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__xnor2_1 _17590_ (.A(_10088_),
    .B(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__or2b_1 _17591_ (.A(_10011_),
    .B_N(_10013_),
    .X(_10157_));
 sky130_fd_sc_hd__a21boi_1 _17592_ (.A1(_09955_),
    .A2(_10014_),
    .B1_N(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__xor2_1 _17593_ (.A(_10156_),
    .B(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__xnor2_1 _17594_ (.A(_10048_),
    .B(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__or2b_1 _17595_ (.A(_10015_),
    .B_N(_10017_),
    .X(_10161_));
 sky130_fd_sc_hd__a21boi_1 _17596_ (.A1(_09918_),
    .A2(_10018_),
    .B1_N(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__xor2_1 _17597_ (.A(_10160_),
    .B(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__xnor2_1 _17598_ (.A(_10039_),
    .B(_10163_),
    .Y(_10164_));
 sky130_fd_sc_hd__and3_1 _17599_ (.A(_10037_),
    .B(_10038_),
    .C(_10164_),
    .X(_10165_));
 sky130_fd_sc_hd__a21o_1 _17600_ (.A1(_10037_),
    .A2(_10038_),
    .B1(_10164_),
    .X(_10166_));
 sky130_fd_sc_hd__or2b_1 _17601_ (.A(_10165_),
    .B_N(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__and2_1 _17602_ (.A(_10023_),
    .B(_10025_),
    .X(_10168_));
 sky130_fd_sc_hd__or2_1 _17603_ (.A(_10023_),
    .B(_10025_),
    .X(_10169_));
 sky130_fd_sc_hd__o21a_1 _17604_ (.A1(_09906_),
    .A2(_10168_),
    .B1(_10169_),
    .X(_10170_));
 sky130_fd_sc_hd__xnor2_2 _17605_ (.A(_10167_),
    .B(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__or2_1 _17606_ (.A(_05203_),
    .B(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__inv_2 _17607_ (.A(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__or2_1 _17608_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_10174_));
 sky130_fd_sc_hd__nand2_1 _17609_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_10175_));
 sky130_fd_sc_hd__a211o_1 _17610_ (.A1(_10174_),
    .A2(_10175_),
    .B1(_10031_),
    .C1(_10033_),
    .X(_10176_));
 sky130_fd_sc_hd__o211ai_2 _17611_ (.A1(_10031_),
    .A2(_10033_),
    .B1(_10174_),
    .C1(_10175_),
    .Y(_10177_));
 sky130_fd_sc_hd__a31o_1 _17612_ (.A1(_09889_),
    .A2(_10176_),
    .A3(_10177_),
    .B1(_09780_),
    .X(_10178_));
 sky130_fd_sc_hd__o22a_1 _17613_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_09817_),
    .B1(_10173_),
    .B2(_10178_),
    .X(_00590_));
 sky130_fd_sc_hd__and2_1 _17614_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_10179_));
 sky130_fd_sc_hd__nor2_1 _17615_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_10180_));
 sky130_fd_sc_hd__a211oi_1 _17616_ (.A1(_10175_),
    .A2(_10177_),
    .B1(_10179_),
    .C1(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__o211a_1 _17617_ (.A1(_10179_),
    .A2(_10180_),
    .B1(_10175_),
    .C1(_10177_),
    .X(_10182_));
 sky130_fd_sc_hd__nand3b_1 _17618_ (.A_N(_10165_),
    .B(_10166_),
    .C(_10026_),
    .Y(_10183_));
 sky130_fd_sc_hd__nor2_1 _17619_ (.A(_09906_),
    .B(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__a21oi_1 _17620_ (.A1(_10169_),
    .A2(_10166_),
    .B1(_10165_),
    .Y(_10185_));
 sky130_fd_sc_hd__a21o_1 _17621_ (.A1(_09912_),
    .A2(_10047_),
    .B1(_10045_),
    .X(_10186_));
 sky130_fd_sc_hd__or2b_1 _17622_ (.A(_10087_),
    .B_N(_10050_),
    .X(_10187_));
 sky130_fd_sc_hd__a21boi_1 _17623_ (.A1(_10053_),
    .A2(_10056_),
    .B1_N(_10054_),
    .Y(_10188_));
 sky130_fd_sc_hd__a21o_1 _17624_ (.A1(_10064_),
    .A2(_10067_),
    .B1(_10188_),
    .X(_10189_));
 sky130_fd_sc_hd__nand3_1 _17625_ (.A(_10064_),
    .B(_10067_),
    .C(_10188_),
    .Y(_10190_));
 sky130_fd_sc_hd__nand2_1 _17626_ (.A(_10189_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__a21oi_1 _17627_ (.A1(_10085_),
    .A2(_10187_),
    .B1(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__and3_1 _17628_ (.A(_10085_),
    .B(_10187_),
    .C(_10191_),
    .X(_10193_));
 sky130_fd_sc_hd__nor2_1 _17629_ (.A(_10192_),
    .B(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__xor2_1 _17630_ (.A(_10042_),
    .B(_10194_),
    .X(_10195_));
 sky130_fd_sc_hd__nor2_1 _17631_ (.A(_10080_),
    .B(_10082_),
    .Y(_10196_));
 sky130_fd_sc_hd__a21o_1 _17632_ (.A1(_10069_),
    .A2(_10083_),
    .B1(_10196_),
    .X(_10197_));
 sky130_fd_sc_hd__nor2_1 _17633_ (.A(_10092_),
    .B(_10107_),
    .Y(_10198_));
 sky130_fd_sc_hd__a21o_1 _17634_ (.A1(_10090_),
    .A2(_10108_),
    .B1(_10198_),
    .X(_10199_));
 sky130_fd_sc_hd__or3_1 _17635_ (.A(_09096_),
    .B(_09480_),
    .C(_09484_),
    .X(_10200_));
 sky130_fd_sc_hd__o22a_1 _17636_ (.A1(_09096_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_09368_),
    .X(_10201_));
 sky130_fd_sc_hd__o21bai_1 _17637_ (.A1(_09368_),
    .A2(_10200_),
    .B1_N(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__nor2_1 _17638_ (.A(_08037_),
    .B(_09704_),
    .Y(_10203_));
 sky130_fd_sc_hd__xnor2_1 _17639_ (.A(_10202_),
    .B(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__or3_1 _17640_ (.A(_08705_),
    .B(_09029_),
    .C(_09165_),
    .X(_10205_));
 sky130_fd_sc_hd__o22a_1 _17641_ (.A1(_09526_),
    .A2(_09029_),
    .B1(_09165_),
    .B2(_09245_),
    .X(_10206_));
 sky130_fd_sc_hd__o21ba_1 _17642_ (.A1(_09391_),
    .A2(_10205_),
    .B1_N(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__nor2_1 _17643_ (.A(_09249_),
    .B(_09359_),
    .Y(_10208_));
 sky130_fd_sc_hd__xnor2_1 _17644_ (.A(_10207_),
    .B(_10208_),
    .Y(_10209_));
 sky130_fd_sc_hd__o31a_1 _17645_ (.A1(_09096_),
    .A2(_09359_),
    .A3(_10060_),
    .B1(_10059_),
    .X(_10210_));
 sky130_fd_sc_hd__nor2_1 _17646_ (.A(_10209_),
    .B(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__and2_1 _17647_ (.A(_10209_),
    .B(_10210_),
    .X(_10212_));
 sky130_fd_sc_hd__nor2_1 _17648_ (.A(_10211_),
    .B(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__xor2_1 _17649_ (.A(_10204_),
    .B(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__a21bo_1 _17650_ (.A1(_10073_),
    .A2(_10077_),
    .B1_N(_10075_),
    .X(_10215_));
 sky130_fd_sc_hd__a21bo_1 _17651_ (.A1(_10095_),
    .A2(_10097_),
    .B1_N(_10093_),
    .X(_10216_));
 sky130_fd_sc_hd__nand2_1 _17652_ (.A(_08445_),
    .B(_08418_),
    .Y(_10217_));
 sky130_fd_sc_hd__xnor2_1 _17653_ (.A(_10074_),
    .B(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__or3_1 _17654_ (.A(_09522_),
    .B(_08425_),
    .C(_10218_),
    .X(_10219_));
 sky130_fd_sc_hd__o21ai_1 _17655_ (.A1(_09522_),
    .A2(_08427_),
    .B1(_10218_),
    .Y(_10220_));
 sky130_fd_sc_hd__and2_1 _17656_ (.A(_10219_),
    .B(_10220_),
    .X(_10221_));
 sky130_fd_sc_hd__and2_1 _17657_ (.A(_10216_),
    .B(_10221_),
    .X(_10222_));
 sky130_fd_sc_hd__or2_1 _17658_ (.A(_10216_),
    .B(_10221_),
    .X(_10223_));
 sky130_fd_sc_hd__and2b_1 _17659_ (.A_N(_10222_),
    .B(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__xnor2_1 _17660_ (.A(_10215_),
    .B(_10224_),
    .Y(_10225_));
 sky130_fd_sc_hd__a21oi_1 _17661_ (.A1(_10071_),
    .A2(_09961_),
    .B1(_10078_),
    .Y(_10226_));
 sky130_fd_sc_hd__a21oi_1 _17662_ (.A1(_10070_),
    .A2(_10079_),
    .B1(_10226_),
    .Y(_10227_));
 sky130_fd_sc_hd__nor2_1 _17663_ (.A(_10225_),
    .B(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__and2_1 _17664_ (.A(_10225_),
    .B(_10227_),
    .X(_10229_));
 sky130_fd_sc_hd__nor2_1 _17665_ (.A(_10228_),
    .B(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__xor2_1 _17666_ (.A(_10214_),
    .B(_10230_),
    .X(_10231_));
 sky130_fd_sc_hd__xnor2_1 _17667_ (.A(_10199_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__xnor2_1 _17668_ (.A(_10197_),
    .B(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__nor2_1 _17669_ (.A(_10103_),
    .B(_10105_),
    .Y(_10234_));
 sky130_fd_sc_hd__a21o_1 _17670_ (.A1(_10098_),
    .A2(_10106_),
    .B1(_10234_),
    .X(_10235_));
 sky130_fd_sc_hd__a21oi_2 _17671_ (.A1(_10112_),
    .A2(_10120_),
    .B1(_10119_),
    .Y(_10236_));
 sky130_fd_sc_hd__or4_1 _17672_ (.A(_08259_),
    .B(_09126_),
    .C(_08493_),
    .D(_08044_),
    .X(_10237_));
 sky130_fd_sc_hd__clkbuf_4 _17673_ (.A(_08044_),
    .X(_10238_));
 sky130_fd_sc_hd__clkbuf_4 _17674_ (.A(_08259_),
    .X(_10239_));
 sky130_fd_sc_hd__o22ai_1 _17675_ (.A1(_09126_),
    .A2(_08493_),
    .B1(_10238_),
    .B2(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__nand2_1 _17676_ (.A(_10237_),
    .B(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__nor2_1 _17677_ (.A(_10094_),
    .B(_08057_),
    .Y(_10242_));
 sky130_fd_sc_hd__xnor2_2 _17678_ (.A(_10241_),
    .B(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__nor2_2 _17679_ (.A(_08802_),
    .B(_09552_),
    .Y(_10244_));
 sky130_fd_sc_hd__xnor2_2 _17680_ (.A(_10099_),
    .B(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__nor2_1 _17681_ (.A(_09276_),
    .B(_09674_),
    .Y(_10246_));
 sky130_fd_sc_hd__xor2_2 _17682_ (.A(_10245_),
    .B(_10246_),
    .X(_10247_));
 sky130_fd_sc_hd__clkbuf_4 _17683_ (.A(_09674_),
    .X(_10248_));
 sky130_fd_sc_hd__nand2_1 _17684_ (.A(_09670_),
    .B(_10099_),
    .Y(_10249_));
 sky130_fd_sc_hd__o31a_1 _17685_ (.A1(_09126_),
    .A2(_10248_),
    .A3(_10100_),
    .B1(_10249_),
    .X(_10250_));
 sky130_fd_sc_hd__xor2_2 _17686_ (.A(_10247_),
    .B(_10250_),
    .X(_10251_));
 sky130_fd_sc_hd__xnor2_2 _17687_ (.A(_10243_),
    .B(_10251_),
    .Y(_10252_));
 sky130_fd_sc_hd__xor2_2 _17688_ (.A(_10236_),
    .B(_10252_),
    .X(_10253_));
 sky130_fd_sc_hd__xor2_2 _17689_ (.A(_10235_),
    .B(_10253_),
    .X(_10254_));
 sky130_fd_sc_hd__nor2_1 _17690_ (.A(_08767_),
    .B(_09693_),
    .Y(_10255_));
 sky130_fd_sc_hd__or2_1 _17691_ (.A(_09980_),
    .B(_10115_),
    .X(_10256_));
 sky130_fd_sc_hd__a22o_1 _17692_ (.A1(_09974_),
    .A2(_10255_),
    .B1(_10256_),
    .B2(_10117_),
    .X(_10257_));
 sky130_fd_sc_hd__a21bo_1 _17693_ (.A1(_10137_),
    .A2(_10141_),
    .B1_N(_10140_),
    .X(_10258_));
 sky130_fd_sc_hd__a21oi_1 _17694_ (.A1(_09292_),
    .A2(_09695_),
    .B1(_08895_),
    .Y(_10259_));
 sky130_fd_sc_hd__xnor2_1 _17695_ (.A(_10255_),
    .B(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__nor2_1 _17696_ (.A(_10110_),
    .B(_09973_),
    .Y(_10261_));
 sky130_fd_sc_hd__xnor2_1 _17697_ (.A(_10260_),
    .B(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__xor2_2 _17698_ (.A(_10258_),
    .B(_10262_),
    .X(_10263_));
 sky130_fd_sc_hd__xor2_2 _17699_ (.A(_10257_),
    .B(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__nor2_1 _17700_ (.A(_09117_),
    .B(_09991_),
    .Y(_10265_));
 sky130_fd_sc_hd__clkbuf_4 _17701_ (.A(_10139_),
    .X(_10266_));
 sky130_fd_sc_hd__a2bb2o_1 _17702_ (.A1_N(_10139_),
    .A2_N(_08873_),
    .B1(_08263_),
    .B2(_10134_),
    .X(_10267_));
 sky130_fd_sc_hd__o21a_1 _17703_ (.A1(_10130_),
    .A2(_10266_),
    .B1(_10267_),
    .X(_10268_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_10265_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__and3_1 _17705_ (.A(_10125_),
    .B(_10133_),
    .C(_10135_),
    .X(_10270_));
 sky130_fd_sc_hd__buf_4 _17706_ (.A(_10270_),
    .X(_10271_));
 sky130_fd_sc_hd__a21oi_2 _17707_ (.A1(_10126_),
    .A2(_10269_),
    .B1(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__xnor2_2 _17708_ (.A(_10264_),
    .B(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__a21oi_1 _17709_ (.A1(_10123_),
    .A2(_10148_),
    .B1(_10145_),
    .Y(_10274_));
 sky130_fd_sc_hd__a21o_1 _17710_ (.A1(_10122_),
    .A2(_10146_),
    .B1(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__xnor2_2 _17711_ (.A(_10273_),
    .B(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__xnor2_2 _17712_ (.A(_10254_),
    .B(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__or2b_1 _17713_ (.A(_10147_),
    .B_N(_10150_),
    .X(_10278_));
 sky130_fd_sc_hd__a21bo_1 _17714_ (.A1(_10109_),
    .A2(_10151_),
    .B1_N(_10278_),
    .X(_10279_));
 sky130_fd_sc_hd__xnor2_1 _17715_ (.A(_10277_),
    .B(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__xnor2_1 _17716_ (.A(_10233_),
    .B(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__nor2_1 _17717_ (.A(_10152_),
    .B(_10154_),
    .Y(_10282_));
 sky130_fd_sc_hd__a21oi_1 _17718_ (.A1(_10088_),
    .A2(_10155_),
    .B1(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__xor2_1 _17719_ (.A(_10281_),
    .B(_10283_),
    .X(_10284_));
 sky130_fd_sc_hd__xnor2_1 _17720_ (.A(_10195_),
    .B(_10284_),
    .Y(_10285_));
 sky130_fd_sc_hd__nor2_1 _17721_ (.A(_10156_),
    .B(_10158_),
    .Y(_10286_));
 sky130_fd_sc_hd__a21oi_1 _17722_ (.A1(_10048_),
    .A2(_10159_),
    .B1(_10286_),
    .Y(_10287_));
 sky130_fd_sc_hd__xor2_1 _17723_ (.A(_10285_),
    .B(_10287_),
    .X(_10288_));
 sky130_fd_sc_hd__xnor2_1 _17724_ (.A(_10186_),
    .B(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__nor2_1 _17725_ (.A(_10160_),
    .B(_10162_),
    .Y(_10290_));
 sky130_fd_sc_hd__a21oi_1 _17726_ (.A1(_10039_),
    .A2(_10163_),
    .B1(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__nor2_1 _17727_ (.A(_10289_),
    .B(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__and2_1 _17728_ (.A(_10289_),
    .B(_10291_),
    .X(_10293_));
 sky130_fd_sc_hd__nor2_1 _17729_ (.A(_10292_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__o21a_1 _17730_ (.A1(_10184_),
    .A2(_10185_),
    .B1(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__or3_1 _17731_ (.A(_10294_),
    .B(_10184_),
    .C(_10185_),
    .X(_10296_));
 sky130_fd_sc_hd__and2b_2 _17732_ (.A_N(_10295_),
    .B(_10296_),
    .X(_10297_));
 sky130_fd_sc_hd__nand2_1 _17733_ (.A(_09812_),
    .B(_10297_),
    .Y(_01438_));
 sky130_fd_sc_hd__o311a_1 _17734_ (.A1(_09812_),
    .A2(_10181_),
    .A3(_10182_),
    .B1(_05414_),
    .C1(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__a21oi_1 _17735_ (.A1(_05268_),
    .A2(_09781_),
    .B1(_01439_),
    .Y(_00591_));
 sky130_fd_sc_hd__nor2_1 _17736_ (.A(_10285_),
    .B(_10287_),
    .Y(_01440_));
 sky130_fd_sc_hd__a21o_1 _17737_ (.A1(_10186_),
    .A2(_10288_),
    .B1(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__a21o_1 _17738_ (.A1(_10042_),
    .A2(_10194_),
    .B1(_10192_),
    .X(_01442_));
 sky130_fd_sc_hd__nand2_1 _17739_ (.A(_10199_),
    .B(_10231_),
    .Y(_01443_));
 sky130_fd_sc_hd__or2b_1 _17740_ (.A(_10232_),
    .B_N(_10197_),
    .X(_01444_));
 sky130_fd_sc_hd__a21o_1 _17741_ (.A1(_10204_),
    .A2(_10213_),
    .B1(_10211_),
    .X(_01445_));
 sky130_fd_sc_hd__o32a_1 _17742_ (.A1(_08331_),
    .A2(_09610_),
    .A3(_10201_),
    .B1(_10200_),
    .B2(_09368_),
    .X(_01446_));
 sky130_fd_sc_hd__inv_2 _17743_ (.A(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _17744_ (.A(_01445_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__or2_1 _17745_ (.A(_01445_),
    .B(_01447_),
    .X(_01449_));
 sky130_fd_sc_hd__nand2_1 _17746_ (.A(_01448_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__a21oi_1 _17747_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__and3_1 _17748_ (.A(_01443_),
    .B(_01444_),
    .C(_01450_),
    .X(_01452_));
 sky130_fd_sc_hd__nor2_1 _17749_ (.A(_01451_),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__xnor2_1 _17750_ (.A(_10189_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__a21o_1 _17751_ (.A1(_10214_),
    .A2(_10230_),
    .B1(_10228_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2_1 _17752_ (.A(_10236_),
    .B(_10252_),
    .Y(_01456_));
 sky130_fd_sc_hd__a21o_1 _17753_ (.A1(_10235_),
    .A2(_10253_),
    .B1(_01456_),
    .X(_01457_));
 sky130_fd_sc_hd__o22a_1 _17754_ (.A1(_09249_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_09096_),
    .X(_01458_));
 sky130_fd_sc_hd__o21ba_1 _17755_ (.A1(_09249_),
    .A2(_10200_),
    .B1_N(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__nand2_1 _17756_ (.A(_09368_),
    .B(_09703_),
    .Y(_01460_));
 sky130_fd_sc_hd__xnor2_1 _17757_ (.A(_01459_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__buf_2 _17758_ (.A(_09522_),
    .X(_01462_));
 sky130_fd_sc_hd__o22a_1 _17759_ (.A1(_01462_),
    .A2(_09029_),
    .B1(_09165_),
    .B2(_09526_),
    .X(_01463_));
 sky130_fd_sc_hd__o21ba_1 _17760_ (.A1(_01462_),
    .A2(_10205_),
    .B1_N(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__nor2_1 _17761_ (.A(_09391_),
    .B(_09359_),
    .Y(_01465_));
 sky130_fd_sc_hd__xnor2_1 _17762_ (.A(_01464_),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__o32a_1 _17763_ (.A1(_09249_),
    .A2(_09359_),
    .A3(_10206_),
    .B1(_10205_),
    .B2(_09391_),
    .X(_01467_));
 sky130_fd_sc_hd__nor2_1 _17764_ (.A(_01466_),
    .B(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__and2_1 _17765_ (.A(_01466_),
    .B(_01467_),
    .X(_01469_));
 sky130_fd_sc_hd__nor2_1 _17766_ (.A(_01468_),
    .B(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__xor2_1 _17767_ (.A(_01461_),
    .B(_01470_),
    .X(_01471_));
 sky130_fd_sc_hd__o21ai_1 _17768_ (.A1(_10074_),
    .A2(_10217_),
    .B1(_10219_),
    .Y(_01472_));
 sky130_fd_sc_hd__a21bo_1 _17769_ (.A1(_10240_),
    .A2(_10242_),
    .B1_N(_10237_),
    .X(_01473_));
 sky130_fd_sc_hd__nand2_2 _17770_ (.A(_05198_),
    .B(_08445_),
    .Y(_01474_));
 sky130_fd_sc_hd__clkbuf_4 _17771_ (.A(_08157_),
    .X(_01475_));
 sky130_fd_sc_hd__clkbuf_4 _17772_ (.A(_08149_),
    .X(_01476_));
 sky130_fd_sc_hd__or4_1 _17773_ (.A(_01474_),
    .B(_08202_),
    .C(_01475_),
    .D(_01476_),
    .X(_01477_));
 sky130_fd_sc_hd__a2bb2o_1 _17774_ (.A1_N(_08202_),
    .A2_N(_01476_),
    .B1(_08417_),
    .B2(_08445_),
    .X(_01478_));
 sky130_fd_sc_hd__nand2_1 _17775_ (.A(_01477_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _17776_ (.A(_07974_),
    .B(_08427_),
    .Y(_01480_));
 sky130_fd_sc_hd__xnor2_1 _17777_ (.A(_01479_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__and2_1 _17778_ (.A(_01473_),
    .B(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__or2_1 _17779_ (.A(_01473_),
    .B(_01481_),
    .X(_01483_));
 sky130_fd_sc_hd__and2b_1 _17780_ (.A_N(_01482_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__xnor2_1 _17781_ (.A(_01472_),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21oi_1 _17782_ (.A1(_10215_),
    .A2(_10224_),
    .B1(_10222_),
    .Y(_01486_));
 sky130_fd_sc_hd__nor2_1 _17783_ (.A(_01485_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__and2_1 _17784_ (.A(_01485_),
    .B(_01486_),
    .X(_01488_));
 sky130_fd_sc_hd__nor2_1 _17785_ (.A(_01487_),
    .B(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__xor2_1 _17786_ (.A(_01471_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__xnor2_1 _17787_ (.A(_01457_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__xnor2_1 _17788_ (.A(_01455_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _17789_ (.A(_10247_),
    .B(_10250_),
    .Y(_01493_));
 sky130_fd_sc_hd__a21o_1 _17790_ (.A1(_10243_),
    .A2(_10251_),
    .B1(_01493_),
    .X(_01494_));
 sky130_fd_sc_hd__and2_1 _17791_ (.A(_10258_),
    .B(_10262_),
    .X(_01495_));
 sky130_fd_sc_hd__a21oi_2 _17792_ (.A1(_10257_),
    .A2(_10263_),
    .B1(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__or4_1 _17793_ (.A(_08188_),
    .B(_09276_),
    .C(_08493_),
    .D(_08044_),
    .X(_01497_));
 sky130_fd_sc_hd__clkbuf_4 _17794_ (.A(_08188_),
    .X(_01498_));
 sky130_fd_sc_hd__o22ai_1 _17795_ (.A1(_09276_),
    .A2(_08493_),
    .B1(_08044_),
    .B2(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_1 _17796_ (.A(_01497_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _17797_ (.A(_10239_),
    .B(_08057_),
    .Y(_01501_));
 sky130_fd_sc_hd__xnor2_2 _17798_ (.A(_01500_),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _17799_ (.A(_09668_),
    .B(_09973_),
    .Y(_01503_));
 sky130_fd_sc_hd__o22a_1 _17800_ (.A1(_09668_),
    .A2(_09552_),
    .B1(_09973_),
    .B2(_08802_),
    .X(_01504_));
 sky130_fd_sc_hd__a21o_1 _17801_ (.A1(_10244_),
    .A2(_01503_),
    .B1(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__nor2_1 _17802_ (.A(_09674_),
    .B(_09417_),
    .Y(_01506_));
 sky130_fd_sc_hd__xor2_2 _17803_ (.A(_01505_),
    .B(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__nand2_1 _17804_ (.A(_10099_),
    .B(_10244_),
    .Y(_01508_));
 sky130_fd_sc_hd__o31a_1 _17805_ (.A1(_09276_),
    .A2(_09674_),
    .A3(_10245_),
    .B1(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__xor2_2 _17806_ (.A(_01507_),
    .B(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__xnor2_2 _17807_ (.A(_01502_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__xor2_2 _17808_ (.A(_01496_),
    .B(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__xor2_2 _17809_ (.A(_01494_),
    .B(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__a21oi_2 _17810_ (.A1(_09292_),
    .A2(_09695_),
    .B1(_08767_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand2_1 _17811_ (.A(_10115_),
    .B(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__o31ai_2 _17812_ (.A1(_10110_),
    .A2(_09973_),
    .A3(_10260_),
    .B1(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__a2bb2o_1 _17813_ (.A1_N(_10130_),
    .A2_N(_10266_),
    .B1(_10265_),
    .B2(_10267_),
    .X(_01517_));
 sky130_fd_sc_hd__a21oi_1 _17814_ (.A1(_09434_),
    .A2(_09988_),
    .B1(_08895_),
    .Y(_01518_));
 sky130_fd_sc_hd__xnor2_1 _17815_ (.A(_01514_),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _17816_ (.A(_09114_),
    .B(_09693_),
    .Y(_01520_));
 sky130_fd_sc_hd__xnor2_1 _17817_ (.A(_01519_),
    .B(_01520_),
    .Y(_01521_));
 sky130_fd_sc_hd__xor2_1 _17818_ (.A(_01517_),
    .B(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__xor2_1 _17819_ (.A(_01516_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__buf_2 _17820_ (.A(_10129_),
    .X(_01524_));
 sky130_fd_sc_hd__and3_1 _17821_ (.A(_08263_),
    .B(_08266_),
    .C(_10134_),
    .X(_01525_));
 sky130_fd_sc_hd__or3b_1 _17822_ (.A(_01524_),
    .B(_01525_),
    .C_N(_10131_),
    .X(_01526_));
 sky130_fd_sc_hd__nor2_1 _17823_ (.A(_09117_),
    .B(_10266_),
    .Y(_01527_));
 sky130_fd_sc_hd__xor2_1 _17824_ (.A(_01526_),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__a21oi_1 _17825_ (.A1(_10126_),
    .A2(_01528_),
    .B1(_10271_),
    .Y(_01529_));
 sky130_fd_sc_hd__xnor2_1 _17826_ (.A(_01523_),
    .B(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__a21oi_1 _17827_ (.A1(_10264_),
    .A2(_10272_),
    .B1(_10271_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _17828_ (.A(_01530_),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _17829_ (.A(_01530_),
    .B(_01531_),
    .Y(_01533_));
 sky130_fd_sc_hd__and2b_1 _17830_ (.A_N(_01532_),
    .B(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__xnor2_2 _17831_ (.A(_01513_),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__or2b_1 _17832_ (.A(_10273_),
    .B_N(_10275_),
    .X(_01536_));
 sky130_fd_sc_hd__a21boi_2 _17833_ (.A1(_10254_),
    .A2(_10276_),
    .B1_N(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__xor2_1 _17834_ (.A(_01535_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__xnor2_1 _17835_ (.A(_01492_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__or2b_1 _17836_ (.A(_10277_),
    .B_N(_10279_),
    .X(_01540_));
 sky130_fd_sc_hd__a21boi_1 _17837_ (.A1(_10233_),
    .A2(_10280_),
    .B1_N(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__xor2_1 _17838_ (.A(_01539_),
    .B(_01541_),
    .X(_01542_));
 sky130_fd_sc_hd__xnor2_1 _17839_ (.A(_01454_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__nor2_1 _17840_ (.A(_10281_),
    .B(_10283_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21oi_1 _17841_ (.A1(_10195_),
    .A2(_10284_),
    .B1(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__xnor2_1 _17842_ (.A(_01543_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__xnor2_1 _17843_ (.A(_01442_),
    .B(_01546_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _17844_ (.A(_01441_),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__and2_1 _17845_ (.A(_01441_),
    .B(_01547_),
    .X(_01549_));
 sky130_fd_sc_hd__nor2_2 _17846_ (.A(_01548_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__nor2_1 _17847_ (.A(_10292_),
    .B(_10295_),
    .Y(_01551_));
 sky130_fd_sc_hd__xnor2_2 _17848_ (.A(_01550_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand2_1 _17849_ (.A(_05532_),
    .B(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_1 _17850_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_01554_));
 sky130_fd_sc_hd__or2_1 _17851_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_01555_));
 sky130_fd_sc_hd__nand2_1 _17852_ (.A(_01554_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__or2_1 _17853_ (.A(_10179_),
    .B(_10181_),
    .X(_01557_));
 sky130_fd_sc_hd__xnor2_1 _17854_ (.A(_01556_),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__a21oi_1 _17855_ (.A1(_09889_),
    .A2(_01558_),
    .B1(_09781_),
    .Y(_01559_));
 sky130_fd_sc_hd__o2bb2a_1 _17856_ (.A1_N(_01553_),
    .A2_N(_01559_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_10036_),
    .X(_00592_));
 sky130_fd_sc_hd__o21bai_1 _17857_ (.A1(_10189_),
    .A2(_01452_),
    .B1_N(_01451_),
    .Y(_01560_));
 sky130_fd_sc_hd__nand2_1 _17858_ (.A(_01457_),
    .B(_01490_),
    .Y(_01561_));
 sky130_fd_sc_hd__or2b_1 _17859_ (.A(_01491_),
    .B_N(_01455_),
    .X(_01562_));
 sky130_fd_sc_hd__a21o_1 _17860_ (.A1(_01461_),
    .A2(_01470_),
    .B1(_01468_),
    .X(_01563_));
 sky130_fd_sc_hd__o22a_1 _17861_ (.A1(_09249_),
    .A2(_10200_),
    .B1(_01458_),
    .B2(_01460_),
    .X(_01564_));
 sky130_fd_sc_hd__inv_2 _17862_ (.A(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _17863_ (.A(_01563_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__or2_1 _17864_ (.A(_01563_),
    .B(_01565_),
    .X(_01567_));
 sky130_fd_sc_hd__nand2_1 _17865_ (.A(_01566_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__a21oi_1 _17866_ (.A1(_01561_),
    .A2(_01562_),
    .B1(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__and3_1 _17867_ (.A(_01561_),
    .B(_01562_),
    .C(_01568_),
    .X(_01570_));
 sky130_fd_sc_hd__nor2_1 _17868_ (.A(_01569_),
    .B(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__xnor2_1 _17869_ (.A(_01448_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__a21o_1 _17870_ (.A1(_01471_),
    .A2(_01489_),
    .B1(_01487_),
    .X(_01573_));
 sky130_fd_sc_hd__nor2_1 _17871_ (.A(_01496_),
    .B(_01511_),
    .Y(_01574_));
 sky130_fd_sc_hd__a21oi_1 _17872_ (.A1(_01494_),
    .A2(_01512_),
    .B1(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__or3_1 _17873_ (.A(_09391_),
    .B(_09351_),
    .C(_09483_),
    .X(_01576_));
 sky130_fd_sc_hd__o22a_1 _17874_ (.A1(_09391_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_09249_),
    .X(_01577_));
 sky130_fd_sc_hd__o21ba_1 _17875_ (.A1(_09249_),
    .A2(_01576_),
    .B1_N(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_09096_),
    .B(_09703_),
    .Y(_01579_));
 sky130_fd_sc_hd__xnor2_1 _17877_ (.A(_01578_),
    .B(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__o22ai_1 _17878_ (.A1(_09661_),
    .A2(_09029_),
    .B1(_09165_),
    .B2(_01462_),
    .Y(_01581_));
 sky130_fd_sc_hd__or2_1 _17879_ (.A(_07974_),
    .B(_09164_),
    .X(_01582_));
 sky130_fd_sc_hd__or3_1 _17880_ (.A(_09522_),
    .B(_09029_),
    .C(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__nand2_1 _17881_ (.A(_01581_),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _17882_ (.A(_09526_),
    .B(_09359_),
    .Y(_01585_));
 sky130_fd_sc_hd__xor2_1 _17883_ (.A(_01584_),
    .B(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__o32a_1 _17884_ (.A1(_09391_),
    .A2(_09359_),
    .A3(_01463_),
    .B1(_10205_),
    .B2(_01462_),
    .X(_01587_));
 sky130_fd_sc_hd__nor2_1 _17885_ (.A(_01586_),
    .B(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__and2_1 _17886_ (.A(_01586_),
    .B(_01587_),
    .X(_01589_));
 sky130_fd_sc_hd__nor2_1 _17887_ (.A(_01588_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__xor2_1 _17888_ (.A(_01580_),
    .B(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__a21bo_1 _17889_ (.A1(_01478_),
    .A2(_01480_),
    .B1_N(_01477_),
    .X(_01592_));
 sky130_fd_sc_hd__a21bo_1 _17890_ (.A1(_01499_),
    .A2(_01501_),
    .B1_N(_01497_),
    .X(_01593_));
 sky130_fd_sc_hd__or4_1 _17891_ (.A(_08259_),
    .B(_08202_),
    .C(_08157_),
    .D(_08149_),
    .X(_01594_));
 sky130_fd_sc_hd__o22ai_1 _17892_ (.A1(_08202_),
    .A2(_01475_),
    .B1(_01476_),
    .B2(_08259_),
    .Y(_01595_));
 sky130_fd_sc_hd__nand2_1 _17893_ (.A(_01594_),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_1 _17894_ (.A(_08275_),
    .B(_08427_),
    .Y(_01597_));
 sky130_fd_sc_hd__xnor2_1 _17895_ (.A(_01596_),
    .B(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__and2_1 _17896_ (.A(_01593_),
    .B(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__or2_1 _17897_ (.A(_01593_),
    .B(_01598_),
    .X(_01600_));
 sky130_fd_sc_hd__and2b_1 _17898_ (.A_N(_01599_),
    .B(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__xnor2_1 _17899_ (.A(_01592_),
    .B(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__a21oi_1 _17900_ (.A1(_01472_),
    .A2(_01484_),
    .B1(_01482_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _17901_ (.A(_01602_),
    .B(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__and2_1 _17902_ (.A(_01602_),
    .B(_01603_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _17903_ (.A(_01604_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__xnor2_1 _17904_ (.A(_01591_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__xor2_1 _17905_ (.A(_01575_),
    .B(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__nand2_1 _17906_ (.A(_01573_),
    .B(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__or2_1 _17907_ (.A(_01573_),
    .B(_01608_),
    .X(_01610_));
 sky130_fd_sc_hd__and2_1 _17908_ (.A(_01609_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__nor2_1 _17909_ (.A(_01507_),
    .B(_01509_),
    .Y(_01612_));
 sky130_fd_sc_hd__a21o_1 _17910_ (.A1(_01502_),
    .A2(_01510_),
    .B1(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__and2_1 _17911_ (.A(_01517_),
    .B(_01521_),
    .X(_01614_));
 sky130_fd_sc_hd__a21oi_1 _17912_ (.A1(_01516_),
    .A2(_01522_),
    .B1(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__a21oi_1 _17913_ (.A1(_08242_),
    .A2(_09129_),
    .B1(_08129_),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _17914_ (.A(_08257_),
    .B(_08044_),
    .Y(_01617_));
 sky130_fd_sc_hd__xnor2_1 _17915_ (.A(_01616_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__or3_1 _17916_ (.A(_01498_),
    .B(_08057_),
    .C(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__buf_2 _17917_ (.A(_08057_),
    .X(_01620_));
 sky130_fd_sc_hd__o21ai_1 _17918_ (.A1(_01498_),
    .A2(_01620_),
    .B1(_01618_),
    .Y(_01621_));
 sky130_fd_sc_hd__and2_1 _17919_ (.A(_01619_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__nor2_1 _17920_ (.A(_08802_),
    .B(_09693_),
    .Y(_01623_));
 sky130_fd_sc_hd__xnor2_1 _17921_ (.A(_01503_),
    .B(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__or2_1 _17922_ (.A(_09103_),
    .B(_09552_),
    .X(_01625_));
 sky130_fd_sc_hd__xnor2_1 _17923_ (.A(_01624_),
    .B(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(_10244_),
    .B(_01503_),
    .Y(_01627_));
 sky130_fd_sc_hd__o31a_1 _17925_ (.A1(_09674_),
    .A2(_09417_),
    .A3(_01504_),
    .B1(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__xor2_1 _17926_ (.A(_01626_),
    .B(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__xnor2_1 _17927_ (.A(_01622_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__xor2_1 _17928_ (.A(_01615_),
    .B(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__xor2_1 _17929_ (.A(_01613_),
    .B(_01631_),
    .X(_01632_));
 sky130_fd_sc_hd__nand2_1 _17930_ (.A(_01514_),
    .B(_01518_),
    .Y(_01633_));
 sky130_fd_sc_hd__o31ai_2 _17931_ (.A1(_10110_),
    .A2(_09693_),
    .A3(_01519_),
    .B1(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__a31o_1 _17932_ (.A1(_10134_),
    .A2(_10131_),
    .A3(_01527_),
    .B1(_01525_),
    .X(_01635_));
 sky130_fd_sc_hd__or3b_1 _17933_ (.A(_08767_),
    .B(_10139_),
    .C_N(_01518_),
    .X(_01636_));
 sky130_fd_sc_hd__a2bb2o_1 _17934_ (.A1_N(_08895_),
    .A2_N(_10139_),
    .B1(_08626_),
    .B2(_09989_),
    .X(_01637_));
 sky130_fd_sc_hd__nor2_1 _17935_ (.A(_10110_),
    .B(_09977_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand3_1 _17936_ (.A(_01636_),
    .B(_01637_),
    .C(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__a21o_1 _17937_ (.A1(_01636_),
    .A2(_01637_),
    .B1(_01638_),
    .X(_01640_));
 sky130_fd_sc_hd__nand3_1 _17938_ (.A(_01635_),
    .B(_01639_),
    .C(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__a21o_1 _17939_ (.A1(_01639_),
    .A2(_01640_),
    .B1(_01635_),
    .X(_01642_));
 sky130_fd_sc_hd__nand3_1 _17940_ (.A(_01634_),
    .B(_01641_),
    .C(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__a21o_1 _17941_ (.A1(_01641_),
    .A2(_01642_),
    .B1(_01634_),
    .X(_01644_));
 sky130_fd_sc_hd__a21boi_2 _17942_ (.A1(_10133_),
    .A2(_10135_),
    .B1_N(_10126_),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_4 _17943_ (.A(_10271_),
    .B(_01645_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand3_2 _17944_ (.A(_01643_),
    .B(_01644_),
    .C(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__a21o_1 _17945_ (.A1(_01643_),
    .A2(_01644_),
    .B1(_01646_),
    .X(_01648_));
 sky130_fd_sc_hd__a21o_1 _17946_ (.A1(_01523_),
    .A2(_01529_),
    .B1(_10271_),
    .X(_01649_));
 sky130_fd_sc_hd__and3_1 _17947_ (.A(_01647_),
    .B(_01648_),
    .C(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__a21o_1 _17948_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_01649_),
    .X(_01651_));
 sky130_fd_sc_hd__and2b_1 _17949_ (.A_N(_01650_),
    .B(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__xnor2_1 _17950_ (.A(_01632_),
    .B(_01652_),
    .Y(_01653_));
 sky130_fd_sc_hd__a21oi_1 _17951_ (.A1(_01513_),
    .A2(_01533_),
    .B1(_01532_),
    .Y(_01654_));
 sky130_fd_sc_hd__xor2_1 _17952_ (.A(_01653_),
    .B(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__xor2_1 _17953_ (.A(_01611_),
    .B(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_1 _17954_ (.A(_01535_),
    .B(_01537_),
    .Y(_01657_));
 sky130_fd_sc_hd__a21oi_1 _17955_ (.A1(_01492_),
    .A2(_01538_),
    .B1(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__xnor2_1 _17956_ (.A(_01656_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__xnor2_1 _17957_ (.A(_01572_),
    .B(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_1 _17958_ (.A(_01539_),
    .B(_01541_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21oi_1 _17959_ (.A1(_01454_),
    .A2(_01542_),
    .B1(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__xnor2_1 _17960_ (.A(_01660_),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__xor2_1 _17961_ (.A(_01560_),
    .B(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__or2b_1 _17962_ (.A(_01546_),
    .B_N(_01442_),
    .X(_01665_));
 sky130_fd_sc_hd__o21a_1 _17963_ (.A1(_01543_),
    .A2(_01545_),
    .B1(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__or2_1 _17964_ (.A(_01664_),
    .B(_01666_),
    .X(_01667_));
 sky130_fd_sc_hd__nand2_1 _17965_ (.A(_01664_),
    .B(_01666_),
    .Y(_01668_));
 sky130_fd_sc_hd__nand2_1 _17966_ (.A(_01667_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__or4bb_1 _17967_ (.A(_10183_),
    .B(_09906_),
    .C_N(_10294_),
    .D_N(_01550_),
    .X(_01670_));
 sky130_fd_sc_hd__or2_1 _17968_ (.A(_01441_),
    .B(_01547_),
    .X(_01671_));
 sky130_fd_sc_hd__a21o_1 _17969_ (.A1(_10292_),
    .A2(_01671_),
    .B1(_01549_),
    .X(_01672_));
 sky130_fd_sc_hd__a31oi_2 _17970_ (.A1(_10294_),
    .A2(_10185_),
    .A3(_01550_),
    .B1(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__and3_1 _17971_ (.A(_01669_),
    .B(_01670_),
    .C(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__and2_1 _17972_ (.A(_01670_),
    .B(_01673_),
    .X(_01675_));
 sky130_fd_sc_hd__or2_1 _17973_ (.A(_01669_),
    .B(_01675_),
    .X(_01676_));
 sky130_fd_sc_hd__or3b_2 _17974_ (.A(_05203_),
    .B(_01674_),
    .C_N(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__nor2_1 _17975_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_01678_));
 sky130_fd_sc_hd__and2_1 _17976_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_01679_));
 sky130_fd_sc_hd__a21boi_2 _17977_ (.A1(_01555_),
    .A2(_01557_),
    .B1_N(_01554_),
    .Y(_01680_));
 sky130_fd_sc_hd__o21ai_1 _17978_ (.A1(_01678_),
    .A2(_01679_),
    .B1(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__o31a_1 _17979_ (.A1(_01678_),
    .A2(_01679_),
    .A3(_01680_),
    .B1(_09889_),
    .X(_01682_));
 sky130_fd_sc_hd__a21oi_1 _17980_ (.A1(_01681_),
    .A2(_01682_),
    .B1(_09780_),
    .Y(_01683_));
 sky130_fd_sc_hd__o2bb2a_1 _17981_ (.A1_N(_01677_),
    .A2_N(_01683_),
    .B1(\rbzero.wall_tracer.trackDistX[4] ),
    .B2(_10036_),
    .X(_00593_));
 sky130_fd_sc_hd__or2_1 _17982_ (.A(_01660_),
    .B(_01662_),
    .X(_01684_));
 sky130_fd_sc_hd__or2b_1 _17983_ (.A(_01663_),
    .B_N(_01560_),
    .X(_01685_));
 sky130_fd_sc_hd__a31o_1 _17984_ (.A1(_01445_),
    .A2(_01447_),
    .A3(_01571_),
    .B1(_01569_),
    .X(_01686_));
 sky130_fd_sc_hd__or2_1 _17985_ (.A(_01575_),
    .B(_01607_),
    .X(_01687_));
 sky130_fd_sc_hd__a21o_1 _17986_ (.A1(_01580_),
    .A2(_01590_),
    .B1(_01588_),
    .X(_01688_));
 sky130_fd_sc_hd__o22a_1 _17987_ (.A1(_09249_),
    .A2(_01576_),
    .B1(_01579_),
    .B2(_01577_),
    .X(_01689_));
 sky130_fd_sc_hd__inv_2 _17988_ (.A(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _17989_ (.A(_01688_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__or2_1 _17990_ (.A(_01688_),
    .B(_01690_),
    .X(_01692_));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(_01691_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__a21oi_1 _17992_ (.A1(_01687_),
    .A2(_01609_),
    .B1(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__and3_1 _17993_ (.A(_01687_),
    .B(_01609_),
    .C(_01693_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_1 _17994_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__xnor2_1 _17995_ (.A(_01566_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__a21o_1 _17996_ (.A1(_01591_),
    .A2(_01606_),
    .B1(_01604_),
    .X(_01698_));
 sky130_fd_sc_hd__nor2_1 _17997_ (.A(_01615_),
    .B(_01630_),
    .Y(_01699_));
 sky130_fd_sc_hd__a21oi_1 _17998_ (.A1(_01613_),
    .A2(_01631_),
    .B1(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__o22a_1 _17999_ (.A1(_09526_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_09391_),
    .X(_01701_));
 sky130_fd_sc_hd__nor2_1 _18000_ (.A(_09526_),
    .B(_01576_),
    .Y(_01702_));
 sky130_fd_sc_hd__or2_1 _18001_ (.A(_01701_),
    .B(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__and2_1 _18002_ (.A(_09249_),
    .B(_09703_),
    .X(_01704_));
 sky130_fd_sc_hd__xnor2_1 _18003_ (.A(_01703_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_1 _18004_ (.A(_08445_),
    .B(_09353_),
    .Y(_01706_));
 sky130_fd_sc_hd__xnor2_1 _18005_ (.A(_01582_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__or3_1 _18006_ (.A(_09522_),
    .B(_09217_),
    .C(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__o21ai_1 _18007_ (.A1(_01462_),
    .A2(_09359_),
    .B1(_01707_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _18008_ (.A(_01708_),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__a21boi_1 _18009_ (.A1(_01581_),
    .A2(_01585_),
    .B1_N(_01583_),
    .Y(_01711_));
 sky130_fd_sc_hd__nor2_1 _18010_ (.A(_01710_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__and2_1 _18011_ (.A(_01710_),
    .B(_01711_),
    .X(_01713_));
 sky130_fd_sc_hd__nor2_1 _18012_ (.A(_01712_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__xor2_1 _18013_ (.A(_01705_),
    .B(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__o31a_1 _18014_ (.A1(_01474_),
    .A2(_08423_),
    .A3(_01596_),
    .B1(_01594_),
    .X(_01716_));
 sky130_fd_sc_hd__nand2_1 _18015_ (.A(_01616_),
    .B(_01617_),
    .Y(_01717_));
 sky130_fd_sc_hd__or4_1 _18016_ (.A(_08259_),
    .B(_08188_),
    .C(_08157_),
    .D(_08149_),
    .X(_01718_));
 sky130_fd_sc_hd__o22ai_1 _18017_ (.A1(_08259_),
    .A2(_08157_),
    .B1(_08149_),
    .B2(_08188_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _18018_ (.A(_01718_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _18019_ (.A(_10094_),
    .B(_08423_),
    .Y(_01721_));
 sky130_fd_sc_hd__xnor2_1 _18020_ (.A(_01720_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__inv_2 _18021_ (.A(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21oi_1 _18022_ (.A1(_01717_),
    .A2(_01619_),
    .B1(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__and3_1 _18023_ (.A(_01717_),
    .B(_01619_),
    .C(_01723_),
    .X(_01725_));
 sky130_fd_sc_hd__or3_1 _18024_ (.A(_01716_),
    .B(_01724_),
    .C(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__o21ai_1 _18025_ (.A1(_01724_),
    .A2(_01725_),
    .B1(_01716_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _18026_ (.A(_01726_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__a21oi_1 _18027_ (.A1(_01592_),
    .A2(_01601_),
    .B1(_01599_),
    .Y(_01729_));
 sky130_fd_sc_hd__xor2_1 _18028_ (.A(_01728_),
    .B(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__xnor2_1 _18029_ (.A(_01715_),
    .B(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__xor2_1 _18030_ (.A(_01700_),
    .B(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__xor2_1 _18031_ (.A(_01698_),
    .B(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__nor2_1 _18032_ (.A(_01626_),
    .B(_01628_),
    .Y(_01734_));
 sky130_fd_sc_hd__a21o_1 _18033_ (.A1(_01622_),
    .A2(_01629_),
    .B1(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__a21bo_1 _18034_ (.A1(_01634_),
    .A2(_01642_),
    .B1_N(_01641_),
    .X(_01736_));
 sky130_fd_sc_hd__buf_2 _18035_ (.A(_08493_),
    .X(_01737_));
 sky130_fd_sc_hd__or4_1 _18036_ (.A(_08242_),
    .B(_01737_),
    .C(_10238_),
    .D(_09552_),
    .X(_01738_));
 sky130_fd_sc_hd__buf_2 _18037_ (.A(_08242_),
    .X(_01739_));
 sky130_fd_sc_hd__o22ai_1 _18038_ (.A1(_01739_),
    .A2(_10238_),
    .B1(_09552_),
    .B2(_01737_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _18039_ (.A(_01738_),
    .B(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _18040_ (.A(_08257_),
    .B(_01620_),
    .Y(_01742_));
 sky130_fd_sc_hd__xnor2_2 _18041_ (.A(_01741_),
    .B(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _18042_ (.A(_09668_),
    .B(_09693_),
    .Y(_01744_));
 sky130_fd_sc_hd__a21oi_2 _18043_ (.A1(_09292_),
    .A2(_09695_),
    .B1(_08802_),
    .Y(_01745_));
 sky130_fd_sc_hd__xnor2_1 _18044_ (.A(_01744_),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _18045_ (.A(_09674_),
    .B(_09973_),
    .Y(_01747_));
 sky130_fd_sc_hd__xor2_1 _18046_ (.A(_01746_),
    .B(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__o2bb2a_1 _18047_ (.A1_N(_01503_),
    .A2_N(_01623_),
    .B1(_01624_),
    .B2(_01625_),
    .X(_01749_));
 sky130_fd_sc_hd__xor2_1 _18048_ (.A(_01748_),
    .B(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__xnor2_1 _18049_ (.A(_01743_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__xnor2_1 _18050_ (.A(_01736_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__xor2_1 _18051_ (.A(_01735_),
    .B(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__nand2_1 _18052_ (.A(_10125_),
    .B(_10136_),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_1 _18053_ (.A(_01636_),
    .B(_01639_),
    .Y(_01755_));
 sky130_fd_sc_hd__a21o_2 _18054_ (.A1(_10131_),
    .A2(_10132_),
    .B1(_01525_),
    .X(_01756_));
 sky130_fd_sc_hd__o22ai_1 _18055_ (.A1(_08895_),
    .A2(_01524_),
    .B1(_10266_),
    .B2(_08767_),
    .Y(_01757_));
 sky130_fd_sc_hd__or4_1 _18056_ (.A(_08895_),
    .B(_08767_),
    .C(_01524_),
    .D(_10139_),
    .X(_01758_));
 sky130_fd_sc_hd__nor2_1 _18057_ (.A(_10110_),
    .B(_09991_),
    .Y(_01759_));
 sky130_fd_sc_hd__nand3_1 _18058_ (.A(_01757_),
    .B(_01758_),
    .C(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__a21o_1 _18059_ (.A1(_01757_),
    .A2(_01758_),
    .B1(_01759_),
    .X(_01761_));
 sky130_fd_sc_hd__nand3_1 _18060_ (.A(_01756_),
    .B(_01760_),
    .C(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__a21o_1 _18061_ (.A1(_01760_),
    .A2(_01761_),
    .B1(_01756_),
    .X(_01763_));
 sky130_fd_sc_hd__nand3_1 _18062_ (.A(_01755_),
    .B(_01762_),
    .C(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__a21o_1 _18063_ (.A1(_01762_),
    .A2(_01763_),
    .B1(_01755_),
    .X(_01765_));
 sky130_fd_sc_hd__and3_1 _18064_ (.A(_01646_),
    .B(_01764_),
    .C(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__a21oi_1 _18065_ (.A1(_01764_),
    .A2(_01765_),
    .B1(_01646_),
    .Y(_01767_));
 sky130_fd_sc_hd__a211o_1 _18066_ (.A1(_01754_),
    .A2(_01647_),
    .B1(_01766_),
    .C1(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__o211ai_2 _18067_ (.A1(_01766_),
    .A2(_01767_),
    .B1(_01754_),
    .C1(_01647_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand3_1 _18068_ (.A(_01753_),
    .B(_01768_),
    .C(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__a21o_1 _18069_ (.A1(_01768_),
    .A2(_01769_),
    .B1(_01753_),
    .X(_01771_));
 sky130_fd_sc_hd__a21o_1 _18070_ (.A1(_01632_),
    .A2(_01651_),
    .B1(_01650_),
    .X(_01772_));
 sky130_fd_sc_hd__nand3_1 _18071_ (.A(_01770_),
    .B(_01771_),
    .C(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21o_1 _18072_ (.A1(_01770_),
    .A2(_01771_),
    .B1(_01772_),
    .X(_01774_));
 sky130_fd_sc_hd__and3_1 _18073_ (.A(_01733_),
    .B(_01773_),
    .C(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__a21oi_1 _18074_ (.A1(_01773_),
    .A2(_01774_),
    .B1(_01733_),
    .Y(_01776_));
 sky130_fd_sc_hd__or2_1 _18075_ (.A(_01775_),
    .B(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__nor2_1 _18076_ (.A(_01653_),
    .B(_01654_),
    .Y(_01778_));
 sky130_fd_sc_hd__a21oi_1 _18077_ (.A1(_01611_),
    .A2(_01655_),
    .B1(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__xor2_1 _18078_ (.A(_01777_),
    .B(_01779_),
    .X(_01780_));
 sky130_fd_sc_hd__xnor2_1 _18079_ (.A(_01697_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2b_1 _18080_ (.A(_01658_),
    .B_N(_01656_),
    .X(_01782_));
 sky130_fd_sc_hd__a21boi_1 _18081_ (.A1(_01572_),
    .A2(_01659_),
    .B1_N(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__xnor2_1 _18082_ (.A(_01781_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__xor2_1 _18083_ (.A(_01686_),
    .B(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__a21oi_1 _18084_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__and3_1 _18085_ (.A(_01684_),
    .B(_01685_),
    .C(_01785_),
    .X(_01787_));
 sky130_fd_sc_hd__nor2_1 _18086_ (.A(_01786_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__inv_2 _18087_ (.A(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__and3_1 _18088_ (.A(_01667_),
    .B(_01676_),
    .C(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__a21oi_1 _18089_ (.A1(_01667_),
    .A2(_01676_),
    .B1(_01789_),
    .Y(_01791_));
 sky130_fd_sc_hd__or3_2 _18090_ (.A(_09807_),
    .B(_01790_),
    .C(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__or2_1 _18091_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_01793_));
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_01794_));
 sky130_fd_sc_hd__o21bai_1 _18093_ (.A1(_01678_),
    .A2(_01680_),
    .B1_N(_01679_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21oi_1 _18094_ (.A1(_01793_),
    .A2(_01794_),
    .B1(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__a31o_1 _18095_ (.A1(_01793_),
    .A2(_01794_),
    .A3(_01795_),
    .B1(_09863_),
    .X(_01797_));
 sky130_fd_sc_hd__o21a_1 _18096_ (.A1(_01796_),
    .A2(_01797_),
    .B1(_09817_),
    .X(_01798_));
 sky130_fd_sc_hd__o2bb2a_1 _18097_ (.A1_N(_01792_),
    .A2_N(_01798_),
    .B1(\rbzero.wall_tracer.trackDistX[5] ),
    .B2(_10036_),
    .X(_00594_));
 sky130_fd_sc_hd__a211o_1 _18098_ (.A1(_01670_),
    .A2(_01673_),
    .B1(_01789_),
    .C1(_01669_),
    .X(_01799_));
 sky130_fd_sc_hd__a21o_1 _18099_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01785_),
    .X(_01800_));
 sky130_fd_sc_hd__a21o_1 _18100_ (.A1(_01667_),
    .A2(_01800_),
    .B1(_01787_),
    .X(_01801_));
 sky130_fd_sc_hd__or2_1 _18101_ (.A(_01781_),
    .B(_01783_),
    .X(_01802_));
 sky130_fd_sc_hd__or2b_1 _18102_ (.A(_01784_),
    .B_N(_01686_),
    .X(_01803_));
 sky130_fd_sc_hd__a31o_1 _18103_ (.A1(_01563_),
    .A2(_01565_),
    .A3(_01696_),
    .B1(_01694_),
    .X(_01804_));
 sky130_fd_sc_hd__or2_1 _18104_ (.A(_01700_),
    .B(_01731_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_1 _18105_ (.A(_01698_),
    .B(_01732_),
    .Y(_01806_));
 sky130_fd_sc_hd__a21o_1 _18106_ (.A1(_01705_),
    .A2(_01714_),
    .B1(_01712_),
    .X(_01807_));
 sky130_fd_sc_hd__inv_2 _18107_ (.A(_01701_),
    .Y(_01808_));
 sky130_fd_sc_hd__a21oi_1 _18108_ (.A1(_01808_),
    .A2(_01704_),
    .B1(_01702_),
    .Y(_01809_));
 sky130_fd_sc_hd__inv_2 _18109_ (.A(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__nand2_1 _18110_ (.A(_01807_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__or2_1 _18111_ (.A(_01807_),
    .B(_01810_),
    .X(_01812_));
 sky130_fd_sc_hd__nand2_1 _18112_ (.A(_01811_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21oi_1 _18113_ (.A1(_01805_),
    .A2(_01806_),
    .B1(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__and3_1 _18114_ (.A(_01805_),
    .B(_01806_),
    .C(_01813_),
    .X(_01815_));
 sky130_fd_sc_hd__nor2_1 _18115_ (.A(_01814_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__xnor2_1 _18116_ (.A(_01691_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _18117_ (.A(_01728_),
    .B(_01729_),
    .Y(_01818_));
 sky130_fd_sc_hd__a21o_1 _18118_ (.A1(_01715_),
    .A2(_01730_),
    .B1(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__and2b_1 _18119_ (.A_N(_01751_),
    .B(_01736_),
    .X(_01820_));
 sky130_fd_sc_hd__a21oi_1 _18120_ (.A1(_01735_),
    .A2(_01752_),
    .B1(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__o22a_1 _18121_ (.A1(_01462_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_09526_),
    .X(_01822_));
 sky130_fd_sc_hd__and4bb_1 _18122_ (.A_N(_01462_),
    .B_N(_09526_),
    .C(_09621_),
    .D(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_01823_));
 sky130_fd_sc_hd__or2_1 _18123_ (.A(_01822_),
    .B(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__and2_1 _18124_ (.A(_09391_),
    .B(_09703_),
    .X(_01825_));
 sky130_fd_sc_hd__xnor2_1 _18125_ (.A(_01824_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _18126_ (.A(_08275_),
    .B(_09165_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _18127_ (.A(_10094_),
    .B(_09027_),
    .Y(_01828_));
 sky130_fd_sc_hd__xnor2_1 _18128_ (.A(_01827_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__or2_1 _18129_ (.A(_07974_),
    .B(_09217_),
    .X(_01830_));
 sky130_fd_sc_hd__xnor2_1 _18130_ (.A(_01829_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__o21a_1 _18131_ (.A1(_01582_),
    .A2(_01706_),
    .B1(_01708_),
    .X(_01832_));
 sky130_fd_sc_hd__or2_1 _18132_ (.A(_01831_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__nand2_1 _18133_ (.A(_01831_),
    .B(_01832_),
    .Y(_01834_));
 sky130_fd_sc_hd__and2_1 _18134_ (.A(_01833_),
    .B(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__nand2_1 _18135_ (.A(_01826_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__or2_1 _18136_ (.A(_01826_),
    .B(_01835_),
    .X(_01837_));
 sky130_fd_sc_hd__and2_1 _18137_ (.A(_01836_),
    .B(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__a21bo_1 _18138_ (.A1(_01719_),
    .A2(_01721_),
    .B1_N(_01718_),
    .X(_01839_));
 sky130_fd_sc_hd__a21bo_1 _18139_ (.A1(_01740_),
    .A2(_01742_),
    .B1_N(_01738_),
    .X(_01840_));
 sky130_fd_sc_hd__nor2_1 _18140_ (.A(_01498_),
    .B(_01475_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_1 _18141_ (.A(_08257_),
    .B(_01476_),
    .Y(_01842_));
 sky130_fd_sc_hd__xnor2_1 _18142_ (.A(_01841_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__or3_1 _18143_ (.A(_10239_),
    .B(_08423_),
    .C(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__o21ai_1 _18144_ (.A1(_10239_),
    .A2(_08423_),
    .B1(_01843_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand2_1 _18145_ (.A(_01844_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__xnor2_2 _18146_ (.A(_01840_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__xnor2_1 _18147_ (.A(_01839_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__o21ba_1 _18148_ (.A1(_01716_),
    .A2(_01725_),
    .B1_N(_01724_),
    .X(_01849_));
 sky130_fd_sc_hd__nor2_1 _18149_ (.A(_01848_),
    .B(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__and2_1 _18150_ (.A(_01848_),
    .B(_01849_),
    .X(_01851_));
 sky130_fd_sc_hd__nor2_1 _18151_ (.A(_01850_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__xnor2_1 _18152_ (.A(_01838_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__xnor2_1 _18153_ (.A(_01821_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__xnor2_1 _18154_ (.A(_01819_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _18155_ (.A(_01748_),
    .B(_01749_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21o_1 _18156_ (.A1(_01743_),
    .A2(_01750_),
    .B1(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__a21bo_1 _18157_ (.A1(_01755_),
    .A2(_01763_),
    .B1_N(_01762_),
    .X(_01858_));
 sky130_fd_sc_hd__or4_2 _18158_ (.A(_08237_),
    .B(_08493_),
    .C(_08044_),
    .D(_09973_),
    .X(_01859_));
 sky130_fd_sc_hd__clkbuf_4 _18159_ (.A(_08237_),
    .X(_01860_));
 sky130_fd_sc_hd__o22ai_1 _18160_ (.A1(_01860_),
    .A2(_10238_),
    .B1(_09973_),
    .B2(_01737_),
    .Y(_01861_));
 sky130_fd_sc_hd__nand2_1 _18161_ (.A(_01859_),
    .B(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__or3_1 _18162_ (.A(_01739_),
    .B(_01620_),
    .C(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__o21ai_1 _18163_ (.A1(_01739_),
    .A2(_01620_),
    .B1(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__and2_1 _18164_ (.A(_01863_),
    .B(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__a21o_1 _18165_ (.A1(_09292_),
    .A2(_09695_),
    .B1(_09668_),
    .X(_01866_));
 sky130_fd_sc_hd__a21oi_1 _18166_ (.A1(_09434_),
    .A2(_09988_),
    .B1(_08802_),
    .Y(_01867_));
 sky130_fd_sc_hd__xnor2_1 _18167_ (.A(_01866_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _18168_ (.A(_09674_),
    .B(_09693_),
    .Y(_01869_));
 sky130_fd_sc_hd__xnor2_1 _18169_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _18170_ (.A(_01744_),
    .B(_01745_),
    .Y(_01871_));
 sky130_fd_sc_hd__o31a_1 _18171_ (.A1(_10248_),
    .A2(_09973_),
    .A3(_01746_),
    .B1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__xor2_1 _18172_ (.A(_01870_),
    .B(_01872_),
    .X(_01873_));
 sky130_fd_sc_hd__xnor2_1 _18173_ (.A(_01865_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__xor2_1 _18174_ (.A(_01858_),
    .B(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__xnor2_1 _18175_ (.A(_01857_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand2_1 _18176_ (.A(_01758_),
    .B(_01760_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand2_1 _18177_ (.A(_08895_),
    .B(_08767_),
    .Y(_01878_));
 sky130_fd_sc_hd__o311a_1 _18178_ (.A1(_08895_),
    .A2(_07916_),
    .A3(_07921_),
    .B1(_10134_),
    .C1(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__nor2_1 _18179_ (.A(_10110_),
    .B(_10266_),
    .Y(_01880_));
 sky130_fd_sc_hd__xor2_1 _18180_ (.A(_01879_),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__xnor2_1 _18181_ (.A(_01756_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__xnor2_1 _18182_ (.A(_01877_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__xnor2_1 _18183_ (.A(_01646_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__o21bai_1 _18184_ (.A1(_10271_),
    .A2(_01766_),
    .B1_N(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__or3b_1 _18185_ (.A(_10271_),
    .B(_01766_),
    .C_N(_01884_),
    .X(_01886_));
 sky130_fd_sc_hd__nand3_1 _18186_ (.A(_01876_),
    .B(_01885_),
    .C(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21o_1 _18187_ (.A1(_01885_),
    .A2(_01886_),
    .B1(_01876_),
    .X(_01888_));
 sky130_fd_sc_hd__a21bo_1 _18188_ (.A1(_01753_),
    .A2(_01769_),
    .B1_N(_01768_),
    .X(_01889_));
 sky130_fd_sc_hd__nand3_1 _18189_ (.A(_01887_),
    .B(_01888_),
    .C(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__a21o_1 _18190_ (.A1(_01887_),
    .A2(_01888_),
    .B1(_01889_),
    .X(_01891_));
 sky130_fd_sc_hd__nand3_1 _18191_ (.A(_01855_),
    .B(_01890_),
    .C(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__a21o_1 _18192_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01855_),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _18193_ (.A(_01892_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__a31o_1 _18194_ (.A1(_01770_),
    .A2(_01771_),
    .A3(_01772_),
    .B1(_01775_),
    .X(_01895_));
 sky130_fd_sc_hd__xnor2_1 _18195_ (.A(_01894_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__xnor2_1 _18196_ (.A(_01817_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__nor2_1 _18197_ (.A(_01777_),
    .B(_01779_),
    .Y(_01898_));
 sky130_fd_sc_hd__a21oi_1 _18198_ (.A1(_01697_),
    .A2(_01780_),
    .B1(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__xnor2_1 _18199_ (.A(_01897_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__xor2_1 _18200_ (.A(_01804_),
    .B(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__a21o_1 _18201_ (.A1(_01802_),
    .A2(_01803_),
    .B1(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__inv_2 _18202_ (.A(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__and3_1 _18203_ (.A(_01802_),
    .B(_01803_),
    .C(_01901_),
    .X(_01904_));
 sky130_fd_sc_hd__or2_1 _18204_ (.A(_01903_),
    .B(_01904_),
    .X(_01905_));
 sky130_fd_sc_hd__a21oi_1 _18205_ (.A1(_01799_),
    .A2(_01801_),
    .B1(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__a31o_1 _18206_ (.A1(_01905_),
    .A2(_01799_),
    .A3(_01801_),
    .B1(_05203_),
    .X(_01907_));
 sky130_fd_sc_hd__or2_1 _18207_ (.A(_01906_),
    .B(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__nor2_1 _18208_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01909_));
 sky130_fd_sc_hd__and2_1 _18209_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .X(_01910_));
 sky130_fd_sc_hd__a21boi_1 _18210_ (.A1(_01793_),
    .A2(_01795_),
    .B1_N(_01794_),
    .Y(_01911_));
 sky130_fd_sc_hd__o21ai_1 _18211_ (.A1(_01909_),
    .A2(_01910_),
    .B1(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__o31a_1 _18212_ (.A1(_01909_),
    .A2(_01910_),
    .A3(_01911_),
    .B1(_05204_),
    .X(_01913_));
 sky130_fd_sc_hd__a21oi_1 _18213_ (.A1(_01912_),
    .A2(_01913_),
    .B1(_09780_),
    .Y(_01914_));
 sky130_fd_sc_hd__o2bb2a_1 _18214_ (.A1_N(_01908_),
    .A2_N(_01914_),
    .B1(\rbzero.wall_tracer.trackDistX[6] ),
    .B2(_10036_),
    .X(_00595_));
 sky130_fd_sc_hd__or2_1 _18215_ (.A(_01897_),
    .B(_01899_),
    .X(_01915_));
 sky130_fd_sc_hd__or2b_1 _18216_ (.A(_01900_),
    .B_N(_01804_),
    .X(_01916_));
 sky130_fd_sc_hd__a31o_1 _18217_ (.A1(_01688_),
    .A2(_01690_),
    .A3(_01816_),
    .B1(_01814_),
    .X(_01917_));
 sky130_fd_sc_hd__or2_1 _18218_ (.A(_01821_),
    .B(_01853_),
    .X(_01918_));
 sky130_fd_sc_hd__or2b_1 _18219_ (.A(_01854_),
    .B_N(_01819_),
    .X(_01919_));
 sky130_fd_sc_hd__inv_2 _18220_ (.A(_01822_),
    .Y(_01920_));
 sky130_fd_sc_hd__a21oi_1 _18221_ (.A1(_01920_),
    .A2(_01825_),
    .B1(_01823_),
    .Y(_01921_));
 sky130_fd_sc_hd__a21o_1 _18222_ (.A1(_01833_),
    .A2(_01836_),
    .B1(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__nand3_1 _18223_ (.A(_01833_),
    .B(_01836_),
    .C(_01921_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand2_1 _18224_ (.A(_01922_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__a21oi_1 _18225_ (.A1(_01918_),
    .A2(_01919_),
    .B1(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__and3_1 _18226_ (.A(_01918_),
    .B(_01919_),
    .C(_01924_),
    .X(_01926_));
 sky130_fd_sc_hd__nor2_1 _18227_ (.A(_01925_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_1 _18228_ (.A(_01811_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__a21o_1 _18229_ (.A1(_01838_),
    .A2(_01852_),
    .B1(_01850_),
    .X(_01929_));
 sky130_fd_sc_hd__or2b_1 _18230_ (.A(_01874_),
    .B_N(_01858_),
    .X(_01930_));
 sky130_fd_sc_hd__or2b_1 _18231_ (.A(_01875_),
    .B_N(_01857_),
    .X(_01931_));
 sky130_fd_sc_hd__nand2_1 _18232_ (.A(_01930_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__o22ai_1 _18233_ (.A1(_09661_),
    .A2(_09480_),
    .B1(_09484_),
    .B2(_01462_),
    .Y(_01933_));
 sky130_fd_sc_hd__or2_2 _18234_ (.A(_09661_),
    .B(_09483_),
    .X(_01934_));
 sky130_fd_sc_hd__or3_1 _18235_ (.A(_01462_),
    .B(_09480_),
    .C(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nand2_1 _18236_ (.A(_01933_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _18237_ (.A(_09526_),
    .B(_09703_),
    .Y(_01937_));
 sky130_fd_sc_hd__xor2_2 _18238_ (.A(_01936_),
    .B(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__nor2_2 _18239_ (.A(_10239_),
    .B(_09027_),
    .Y(_01939_));
 sky130_fd_sc_hd__nor2_1 _18240_ (.A(_10094_),
    .B(_09162_),
    .Y(_01940_));
 sky130_fd_sc_hd__xnor2_2 _18241_ (.A(_01939_),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__or2_1 _18242_ (.A(_08275_),
    .B(_09217_),
    .X(_01942_));
 sky130_fd_sc_hd__xnor2_1 _18243_ (.A(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _18244_ (.A(_01827_),
    .B(_01828_),
    .Y(_01944_));
 sky130_fd_sc_hd__o31a_1 _18245_ (.A1(_09661_),
    .A2(_09359_),
    .A3(_01829_),
    .B1(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__or2_1 _18246_ (.A(_01943_),
    .B(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__nand2_1 _18247_ (.A(_01943_),
    .B(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__and2_1 _18248_ (.A(_01946_),
    .B(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__nand2_1 _18249_ (.A(_01938_),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__or2_1 _18250_ (.A(_01938_),
    .B(_01948_),
    .X(_01950_));
 sky130_fd_sc_hd__and2_1 _18251_ (.A(_01949_),
    .B(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__a21bo_1 _18252_ (.A1(_01841_),
    .A2(_01842_),
    .B1_N(_01844_),
    .X(_01952_));
 sky130_fd_sc_hd__nand2_1 _18253_ (.A(_01859_),
    .B(_01863_),
    .Y(_01953_));
 sky130_fd_sc_hd__or4_1 _18254_ (.A(_08257_),
    .B(_08242_),
    .C(_01475_),
    .D(_01476_),
    .X(_01954_));
 sky130_fd_sc_hd__o22ai_1 _18255_ (.A1(_08257_),
    .A2(_01475_),
    .B1(_01476_),
    .B2(_01739_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _18256_ (.A(_01954_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__nor2_1 _18257_ (.A(_01498_),
    .B(_08423_),
    .Y(_01957_));
 sky130_fd_sc_hd__xor2_1 _18258_ (.A(_01956_),
    .B(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__xnor2_1 _18259_ (.A(_01953_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__xnor2_1 _18260_ (.A(_01952_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__and2b_1 _18261_ (.A_N(_01846_),
    .B(_01840_),
    .X(_01961_));
 sky130_fd_sc_hd__a21oi_2 _18262_ (.A1(_01839_),
    .A2(_01847_),
    .B1(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__xor2_1 _18263_ (.A(_01960_),
    .B(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__xnor2_1 _18264_ (.A(_01951_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__xor2_1 _18265_ (.A(_01932_),
    .B(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__xnor2_2 _18266_ (.A(_01929_),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__or3_1 _18267_ (.A(_08895_),
    .B(_08767_),
    .C(_01524_),
    .X(_01967_));
 sky130_fd_sc_hd__a21bo_1 _18268_ (.A1(_01879_),
    .A2(_01880_),
    .B1_N(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__nor2_1 _18269_ (.A(_10110_),
    .B(_01524_),
    .Y(_01969_));
 sky130_fd_sc_hd__mux2_2 _18270_ (.A0(_01969_),
    .A1(_10110_),
    .S(_01879_),
    .X(_01970_));
 sky130_fd_sc_hd__xnor2_4 _18271_ (.A(_01756_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xnor2_1 _18272_ (.A(_01968_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__xnor2_1 _18273_ (.A(_01646_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__a21oi_1 _18274_ (.A1(_01646_),
    .A2(_01883_),
    .B1(_10271_),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_1 _18275_ (.A(_01973_),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__and2_1 _18276_ (.A(_01973_),
    .B(_01974_),
    .X(_01976_));
 sky130_fd_sc_hd__nor2_1 _18277_ (.A(_01975_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _18278_ (.A(_01870_),
    .B(_01872_),
    .Y(_01978_));
 sky130_fd_sc_hd__a21o_1 _18279_ (.A1(_01865_),
    .A2(_01873_),
    .B1(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__and2b_1 _18280_ (.A_N(_01882_),
    .B(_01877_),
    .X(_01980_));
 sky130_fd_sc_hd__a21o_1 _18281_ (.A1(_01756_),
    .A2(_01881_),
    .B1(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__nor2_1 _18282_ (.A(_01737_),
    .B(_09693_),
    .Y(_01982_));
 sky130_fd_sc_hd__nor2_1 _18283_ (.A(_09141_),
    .B(_10238_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_1 _18284_ (.A(_01982_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__or3_1 _18285_ (.A(_01860_),
    .B(_01620_),
    .C(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__o21ai_1 _18286_ (.A1(_01860_),
    .A2(_01620_),
    .B1(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__and2_1 _18287_ (.A(_01985_),
    .B(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__nor2_1 _18288_ (.A(_09668_),
    .B(_09991_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor2_1 _18289_ (.A(_08802_),
    .B(_10139_),
    .Y(_01989_));
 sky130_fd_sc_hd__xnor2_1 _18290_ (.A(_01988_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _18291_ (.A(_10248_),
    .B(_09977_),
    .Y(_01991_));
 sky130_fd_sc_hd__xor2_1 _18292_ (.A(_01990_),
    .B(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__a22oi_2 _18293_ (.A1(_01745_),
    .A2(_01988_),
    .B1(_01868_),
    .B2(_01869_),
    .Y(_01993_));
 sky130_fd_sc_hd__xor2_1 _18294_ (.A(_01992_),
    .B(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__xnor2_1 _18295_ (.A(_01987_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__xor2_1 _18296_ (.A(_01981_),
    .B(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__xnor2_1 _18297_ (.A(_01979_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__xnor2_2 _18298_ (.A(_01977_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__and2_1 _18299_ (.A(_01885_),
    .B(_01887_),
    .X(_01999_));
 sky130_fd_sc_hd__xor2_2 _18300_ (.A(_01998_),
    .B(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__xnor2_2 _18301_ (.A(_01966_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__and2_1 _18302_ (.A(_01890_),
    .B(_01892_),
    .X(_02002_));
 sky130_fd_sc_hd__nor2_1 _18303_ (.A(_02001_),
    .B(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _18304_ (.A(_02001_),
    .B(_02002_),
    .Y(_02004_));
 sky130_fd_sc_hd__and2b_1 _18305_ (.A_N(_02003_),
    .B(_02004_),
    .X(_02005_));
 sky130_fd_sc_hd__xnor2_1 _18306_ (.A(_01928_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__and3_1 _18307_ (.A(_01892_),
    .B(_01893_),
    .C(_01895_),
    .X(_02007_));
 sky130_fd_sc_hd__a21oi_1 _18308_ (.A1(_01817_),
    .A2(_01896_),
    .B1(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__xnor2_1 _18309_ (.A(_02006_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__xor2_1 _18310_ (.A(_01917_),
    .B(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__and3_1 _18311_ (.A(_01915_),
    .B(_01916_),
    .C(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__a21o_1 _18312_ (.A1(_01915_),
    .A2(_01916_),
    .B1(_02010_),
    .X(_02012_));
 sky130_fd_sc_hd__or2b_1 _18313_ (.A(_02011_),
    .B_N(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__nor2_1 _18314_ (.A(_01903_),
    .B(_01906_),
    .Y(_02014_));
 sky130_fd_sc_hd__xnor2_1 _18315_ (.A(_02013_),
    .B(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__or2_1 _18316_ (.A(_09889_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__or2_1 _18317_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .X(_02017_));
 sky130_fd_sc_hd__nand2_1 _18318_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_02018_));
 sky130_fd_sc_hd__o21bai_1 _18319_ (.A1(_01909_),
    .A2(_01911_),
    .B1_N(_01910_),
    .Y(_02019_));
 sky130_fd_sc_hd__a21oi_1 _18320_ (.A1(_02017_),
    .A2(_02018_),
    .B1(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__a31o_1 _18321_ (.A1(_02017_),
    .A2(_02018_),
    .A3(_02019_),
    .B1(_05531_),
    .X(_02021_));
 sky130_fd_sc_hd__o21a_1 _18322_ (.A1(_02020_),
    .A2(_02021_),
    .B1(_09817_),
    .X(_02022_));
 sky130_fd_sc_hd__o2bb2a_1 _18323_ (.A1_N(_02016_),
    .A2_N(_02022_),
    .B1(\rbzero.wall_tracer.trackDistX[7] ),
    .B2(_10036_),
    .X(_00596_));
 sky130_fd_sc_hd__a21o_1 _18324_ (.A1(_01902_),
    .A2(_02012_),
    .B1(_02011_),
    .X(_02023_));
 sky130_fd_sc_hd__and2_1 _18325_ (.A(_01801_),
    .B(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__or2_1 _18326_ (.A(_01905_),
    .B(_02013_),
    .X(_02025_));
 sky130_fd_sc_hd__nand2_1 _18327_ (.A(_10134_),
    .B(_01878_),
    .Y(_02026_));
 sky130_fd_sc_hd__o21a_1 _18328_ (.A1(_10110_),
    .A2(_02026_),
    .B1(_01967_),
    .X(_02027_));
 sky130_fd_sc_hd__xor2_1 _18329_ (.A(_01971_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__xnor2_1 _18330_ (.A(_01646_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__a21o_1 _18331_ (.A1(_01646_),
    .A2(_01972_),
    .B1(_10271_),
    .X(_02030_));
 sky130_fd_sc_hd__and2b_1 _18332_ (.A_N(_02029_),
    .B(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__and2b_1 _18333_ (.A_N(_02030_),
    .B(_02029_),
    .X(_02032_));
 sky130_fd_sc_hd__nor2_1 _18334_ (.A(_02031_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _18335_ (.A(_01992_),
    .B(_01993_),
    .Y(_02034_));
 sky130_fd_sc_hd__a21o_1 _18336_ (.A1(_01987_),
    .A2(_01994_),
    .B1(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__nand2_1 _18337_ (.A(_01756_),
    .B(_01970_),
    .Y(_02036_));
 sky130_fd_sc_hd__or2b_1 _18338_ (.A(_01971_),
    .B_N(_01968_),
    .X(_02037_));
 sky130_fd_sc_hd__nand2_1 _18339_ (.A(_02036_),
    .B(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__or4_1 _18340_ (.A(_01737_),
    .B(_10238_),
    .C(_09294_),
    .D(_09977_),
    .X(_02039_));
 sky130_fd_sc_hd__o22ai_1 _18341_ (.A1(_10238_),
    .A2(_09294_),
    .B1(_09977_),
    .B2(_01737_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _18342_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__or3_1 _18343_ (.A(_09141_),
    .B(_01620_),
    .C(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__o21ai_1 _18344_ (.A1(_09141_),
    .A2(_01620_),
    .B1(_02041_),
    .Y(_02043_));
 sky130_fd_sc_hd__and2_1 _18345_ (.A(_02042_),
    .B(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__or3_2 _18346_ (.A(_08802_),
    .B(_09668_),
    .C(_01524_),
    .X(_02045_));
 sky130_fd_sc_hd__o22a_1 _18347_ (.A1(_08802_),
    .A2(_01524_),
    .B1(_10139_),
    .B2(_09668_),
    .X(_02046_));
 sky130_fd_sc_hd__o21ba_1 _18348_ (.A1(_10266_),
    .A2(_02045_),
    .B1_N(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__nor2_1 _18349_ (.A(_10248_),
    .B(_09991_),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_1 _18350_ (.A(_02047_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__nand2_1 _18351_ (.A(_01988_),
    .B(_01989_),
    .Y(_02050_));
 sky130_fd_sc_hd__o31a_1 _18352_ (.A1(_10248_),
    .A2(_09977_),
    .A3(_01990_),
    .B1(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__xor2_1 _18353_ (.A(_02049_),
    .B(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__xor2_1 _18354_ (.A(_02044_),
    .B(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__xnor2_1 _18355_ (.A(_02038_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__xnor2_1 _18356_ (.A(_02035_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__xnor2_1 _18357_ (.A(_02033_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__a21oi_1 _18358_ (.A1(_01977_),
    .A2(_01997_),
    .B1(_01975_),
    .Y(_02057_));
 sky130_fd_sc_hd__nor2_1 _18359_ (.A(_02056_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__and2_1 _18360_ (.A(_02056_),
    .B(_02057_),
    .X(_02059_));
 sky130_fd_sc_hd__nor2_1 _18361_ (.A(_02058_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__nor2_1 _18362_ (.A(_01960_),
    .B(_01962_),
    .Y(_02061_));
 sky130_fd_sc_hd__a21o_1 _18363_ (.A1(_01951_),
    .A2(_01963_),
    .B1(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__or2b_1 _18364_ (.A(_01995_),
    .B_N(_01981_),
    .X(_02063_));
 sky130_fd_sc_hd__or2b_1 _18365_ (.A(_01996_),
    .B_N(_01979_),
    .X(_02064_));
 sky130_fd_sc_hd__nand2_1 _18366_ (.A(_02063_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor3_1 _18367_ (.A(_01474_),
    .B(_09350_),
    .C(_01934_),
    .Y(_02066_));
 sky130_fd_sc_hd__o21a_1 _18368_ (.A1(_01474_),
    .A2(_09350_),
    .B1(_01934_),
    .X(_02067_));
 sky130_fd_sc_hd__nor2_1 _18369_ (.A(_02066_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _18370_ (.A(_01462_),
    .B(_09703_),
    .Y(_02069_));
 sky130_fd_sc_hd__xnor2_1 _18371_ (.A(_02068_),
    .B(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _18372_ (.A(_01498_),
    .B(_09162_),
    .Y(_02071_));
 sky130_fd_sc_hd__o22a_1 _18373_ (.A1(_01498_),
    .A2(_09027_),
    .B1(_09162_),
    .B2(_10239_),
    .X(_02072_));
 sky130_fd_sc_hd__a21o_1 _18374_ (.A1(_01939_),
    .A2(_02071_),
    .B1(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__nor2_1 _18375_ (.A(_10094_),
    .B(_09215_),
    .Y(_02074_));
 sky130_fd_sc_hd__xor2_1 _18376_ (.A(_02073_),
    .B(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__nand2_1 _18377_ (.A(_01939_),
    .B(_01940_),
    .Y(_02076_));
 sky130_fd_sc_hd__o31a_1 _18378_ (.A1(_01474_),
    .A2(_09215_),
    .A3(_01941_),
    .B1(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__or2_1 _18379_ (.A(_02075_),
    .B(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__nand2_1 _18380_ (.A(_02075_),
    .B(_02077_),
    .Y(_02079_));
 sky130_fd_sc_hd__and2_1 _18381_ (.A(_02078_),
    .B(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(_02070_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__or2_1 _18383_ (.A(_02070_),
    .B(_02080_),
    .X(_02082_));
 sky130_fd_sc_hd__and2_1 _18384_ (.A(_02081_),
    .B(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__a21bo_1 _18385_ (.A1(_01955_),
    .A2(_01957_),
    .B1_N(_01954_),
    .X(_02084_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(_01982_),
    .B(_01983_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _18387_ (.A(_02085_),
    .B(_01985_),
    .Y(_02086_));
 sky130_fd_sc_hd__or4_1 _18388_ (.A(_01739_),
    .B(_01860_),
    .C(_01475_),
    .D(_01476_),
    .X(_02087_));
 sky130_fd_sc_hd__o22ai_1 _18389_ (.A1(_01739_),
    .A2(_01475_),
    .B1(_01476_),
    .B2(_01860_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_1 _18390_ (.A(_02087_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__nor2_1 _18391_ (.A(_08257_),
    .B(_08423_),
    .Y(_02090_));
 sky130_fd_sc_hd__xor2_1 _18392_ (.A(_02089_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_1 _18393_ (.A(_02086_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__xnor2_1 _18394_ (.A(_02084_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__a21oi_1 _18395_ (.A1(_01859_),
    .A2(_01863_),
    .B1(_01958_),
    .Y(_02094_));
 sky130_fd_sc_hd__a21oi_1 _18396_ (.A1(_01952_),
    .A2(_01959_),
    .B1(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _18397_ (.A(_02093_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_1 _18398_ (.A(_02093_),
    .B(_02095_),
    .Y(_02097_));
 sky130_fd_sc_hd__and2b_1 _18399_ (.A_N(_02096_),
    .B(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__xnor2_1 _18400_ (.A(_02083_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__xor2_1 _18401_ (.A(_02065_),
    .B(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__xnor2_2 _18402_ (.A(_02062_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__xnor2_2 _18403_ (.A(_02060_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _18404_ (.A(_01998_),
    .B(_01999_),
    .Y(_02103_));
 sky130_fd_sc_hd__a21oi_2 _18405_ (.A1(_01966_),
    .A2(_02000_),
    .B1(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__xor2_2 _18406_ (.A(_02102_),
    .B(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__or2b_1 _18407_ (.A(_01964_),
    .B_N(_01932_),
    .X(_02106_));
 sky130_fd_sc_hd__or2b_1 _18408_ (.A(_01965_),
    .B_N(_01929_),
    .X(_02107_));
 sky130_fd_sc_hd__o21a_2 _18409_ (.A1(_01936_),
    .A2(_01937_),
    .B1(_01935_),
    .X(_02108_));
 sky130_fd_sc_hd__a21oi_4 _18410_ (.A1(_01946_),
    .A2(_01949_),
    .B1(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__and3_1 _18411_ (.A(_01946_),
    .B(_01949_),
    .C(_02108_),
    .X(_02110_));
 sky130_fd_sc_hd__or2_1 _18412_ (.A(_02109_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__a21o_1 _18413_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__nand3_1 _18414_ (.A(_02106_),
    .B(_02107_),
    .C(_02111_),
    .Y(_02113_));
 sky130_fd_sc_hd__and2_1 _18415_ (.A(_02112_),
    .B(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__xnor2_1 _18416_ (.A(_01922_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__xnor2_2 _18417_ (.A(_02105_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__a21oi_1 _18418_ (.A1(_01928_),
    .A2(_02004_),
    .B1(_02003_),
    .Y(_02117_));
 sky130_fd_sc_hd__xnor2_1 _18419_ (.A(_02116_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__a31oi_1 _18420_ (.A1(_01807_),
    .A2(_01810_),
    .A3(_01927_),
    .B1(_01925_),
    .Y(_02119_));
 sky130_fd_sc_hd__or2_1 _18421_ (.A(_02118_),
    .B(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__nand2_1 _18422_ (.A(_02118_),
    .B(_02119_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _18423_ (.A(_02120_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__or2b_1 _18424_ (.A(_02009_),
    .B_N(_01917_),
    .X(_02123_));
 sky130_fd_sc_hd__o21a_1 _18425_ (.A1(_02006_),
    .A2(_02008_),
    .B1(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__or2_2 _18426_ (.A(_02122_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__nand2_1 _18427_ (.A(_02122_),
    .B(_02124_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_1 _18428_ (.A(_02125_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__a221o_4 _18429_ (.A1(_01799_),
    .A2(_02024_),
    .B1(_02025_),
    .B2(_02023_),
    .C1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__a22o_1 _18430_ (.A1(_01799_),
    .A2(_02024_),
    .B1(_02025_),
    .B2(_02023_),
    .X(_02129_));
 sky130_fd_sc_hd__a21oi_2 _18431_ (.A1(_02127_),
    .A2(_02129_),
    .B1(_09807_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _18432_ (.A(_02128_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__nor2_1 _18433_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_02132_));
 sky130_fd_sc_hd__and2_1 _18434_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_02133_));
 sky130_fd_sc_hd__a21boi_1 _18435_ (.A1(_02017_),
    .A2(_02019_),
    .B1_N(_02018_),
    .Y(_02134_));
 sky130_fd_sc_hd__o21ai_1 _18436_ (.A1(_02132_),
    .A2(_02133_),
    .B1(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__o31a_1 _18437_ (.A1(_02132_),
    .A2(_02133_),
    .A3(_02134_),
    .B1(_05204_),
    .X(_02136_));
 sky130_fd_sc_hd__a21oi_1 _18438_ (.A1(_02135_),
    .A2(_02136_),
    .B1(_09780_),
    .Y(_02137_));
 sky130_fd_sc_hd__o2bb2a_1 _18439_ (.A1_N(_02131_),
    .A2_N(_02137_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_10036_),
    .X(_00597_));
 sky130_fd_sc_hd__or2_1 _18440_ (.A(_02116_),
    .B(_02117_),
    .X(_02138_));
 sky130_fd_sc_hd__and2b_1 _18441_ (.A_N(_02028_),
    .B(_01645_),
    .X(_02139_));
 sky130_fd_sc_hd__nand2_1 _18442_ (.A(_10271_),
    .B(_02028_),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2b_1 _18443_ (.A(_02139_),
    .B_N(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_1 _18444_ (.A(_02049_),
    .B(_02051_),
    .Y(_02142_));
 sky130_fd_sc_hd__a21o_1 _18445_ (.A1(_02044_),
    .A2(_02052_),
    .B1(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__o21ai_4 _18446_ (.A1(_01971_),
    .A2(_02027_),
    .B1(_02036_),
    .Y(_02144_));
 sky130_fd_sc_hd__or4_1 _18447_ (.A(_01737_),
    .B(_10238_),
    .C(_09292_),
    .D(_09991_),
    .X(_02145_));
 sky130_fd_sc_hd__o22ai_1 _18448_ (.A1(_10238_),
    .A2(_09292_),
    .B1(_09991_),
    .B2(_01737_),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_1 _18449_ (.A(_02145_),
    .B(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__nor2_1 _18450_ (.A(_08356_),
    .B(_09138_),
    .Y(_02148_));
 sky130_fd_sc_hd__xor2_2 _18451_ (.A(_02147_),
    .B(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__a21oi_1 _18452_ (.A1(_08802_),
    .A2(_09668_),
    .B1(_01524_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(_02045_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _18454_ (.A(_10248_),
    .B(_10266_),
    .Y(_02152_));
 sky130_fd_sc_hd__xor2_1 _18455_ (.A(_02151_),
    .B(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__o32a_1 _18456_ (.A1(_10248_),
    .A2(_09991_),
    .A3(_02046_),
    .B1(_02045_),
    .B2(_10266_),
    .X(_02154_));
 sky130_fd_sc_hd__nor2_1 _18457_ (.A(_02153_),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__and2_1 _18458_ (.A(_02153_),
    .B(_02154_),
    .X(_02156_));
 sky130_fd_sc_hd__nor2_1 _18459_ (.A(_02155_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_1 _18460_ (.A(_02149_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__xnor2_1 _18461_ (.A(_02144_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__xnor2_1 _18462_ (.A(_02143_),
    .B(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hd__xnor2_1 _18463_ (.A(_02141_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__a21oi_1 _18464_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_02031_),
    .Y(_02162_));
 sky130_fd_sc_hd__xor2_1 _18465_ (.A(_02161_),
    .B(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__a21o_1 _18466_ (.A1(_02083_),
    .A2(_02097_),
    .B1(_02096_),
    .X(_02164_));
 sky130_fd_sc_hd__or2b_1 _18467_ (.A(_02054_),
    .B_N(_02035_),
    .X(_02165_));
 sky130_fd_sc_hd__a21bo_1 _18468_ (.A1(_02038_),
    .A2(_02053_),
    .B1_N(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__nor2_1 _18469_ (.A(_10094_),
    .B(_09350_),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _18470_ (.A(_08275_),
    .B(_09484_),
    .Y(_02168_));
 sky130_fd_sc_hd__xnor2_1 _18471_ (.A(_02167_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__and2_1 _18472_ (.A(_09661_),
    .B(_09611_),
    .X(_02170_));
 sky130_fd_sc_hd__xnor2_1 _18473_ (.A(_02169_),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _18474_ (.A(_08257_),
    .B(_09027_),
    .Y(_02172_));
 sky130_fd_sc_hd__xnor2_1 _18475_ (.A(_02071_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__or3_1 _18476_ (.A(_10239_),
    .B(_09215_),
    .C(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__o21ai_1 _18477_ (.A1(_10239_),
    .A2(_09215_),
    .B1(_02173_),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _18478_ (.A(_02174_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nand2_1 _18479_ (.A(_01939_),
    .B(_02071_),
    .Y(_02177_));
 sky130_fd_sc_hd__o31a_1 _18480_ (.A1(_10094_),
    .A2(_09215_),
    .A3(_02072_),
    .B1(_02177_),
    .X(_02178_));
 sky130_fd_sc_hd__or2_1 _18481_ (.A(_02176_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__nand2_1 _18482_ (.A(_02176_),
    .B(_02178_),
    .Y(_02180_));
 sky130_fd_sc_hd__and2_1 _18483_ (.A(_02179_),
    .B(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__nand2_1 _18484_ (.A(_02171_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_1 _18485_ (.A(_02171_),
    .B(_02181_),
    .X(_02183_));
 sky130_fd_sc_hd__and2_1 _18486_ (.A(_02182_),
    .B(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__a21bo_1 _18487_ (.A1(_02088_),
    .A2(_02090_),
    .B1_N(_02087_),
    .X(_02185_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(_02039_),
    .B(_02042_),
    .Y(_02186_));
 sky130_fd_sc_hd__or4_1 _18489_ (.A(_01860_),
    .B(_09141_),
    .C(_01475_),
    .D(_01476_),
    .X(_02187_));
 sky130_fd_sc_hd__o22ai_1 _18490_ (.A1(_01860_),
    .A2(_01475_),
    .B1(_01476_),
    .B2(_09141_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _18491_ (.A(_02187_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _18492_ (.A(_01739_),
    .B(_08423_),
    .Y(_02190_));
 sky130_fd_sc_hd__xor2_1 _18493_ (.A(_02189_),
    .B(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__xor2_1 _18494_ (.A(_02186_),
    .B(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__xor2_1 _18495_ (.A(_02185_),
    .B(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__a21oi_1 _18496_ (.A1(_02085_),
    .A2(_01985_),
    .B1(_02091_),
    .Y(_02194_));
 sky130_fd_sc_hd__a21oi_1 _18497_ (.A1(_02084_),
    .A2(_02092_),
    .B1(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__xor2_1 _18498_ (.A(_02193_),
    .B(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__xor2_1 _18499_ (.A(_02184_),
    .B(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__xnor2_1 _18500_ (.A(_02166_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__xnor2_1 _18501_ (.A(_02164_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _18502_ (.A(_02163_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__a21oi_1 _18503_ (.A1(_02060_),
    .A2(_02101_),
    .B1(_02058_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _18504_ (.A(_02200_),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__and2_1 _18505_ (.A(_02200_),
    .B(_02201_),
    .X(_02203_));
 sky130_fd_sc_hd__nor2_1 _18506_ (.A(_02202_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__or2b_1 _18507_ (.A(_02099_),
    .B_N(_02065_),
    .X(_02205_));
 sky130_fd_sc_hd__or2b_1 _18508_ (.A(_02100_),
    .B_N(_02062_),
    .X(_02206_));
 sky130_fd_sc_hd__o21ba_1 _18509_ (.A1(_02067_),
    .A2(_02069_),
    .B1_N(_02066_),
    .X(_02207_));
 sky130_fd_sc_hd__a21o_1 _18510_ (.A1(_02078_),
    .A2(_02081_),
    .B1(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__nand3_1 _18511_ (.A(_02078_),
    .B(_02081_),
    .C(_02207_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _18512_ (.A(_02208_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__a21oi_1 _18513_ (.A1(_02205_),
    .A2(_02206_),
    .B1(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__and3_1 _18514_ (.A(_02205_),
    .B(_02206_),
    .C(_02210_),
    .X(_02212_));
 sky130_fd_sc_hd__nor2_1 _18515_ (.A(_02211_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__xor2_2 _18516_ (.A(_02109_),
    .B(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__xnor2_2 _18517_ (.A(_02204_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _18518_ (.A(_02102_),
    .B(_02104_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21oi_1 _18519_ (.A1(_02105_),
    .A2(_02115_),
    .B1(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__xnor2_2 _18520_ (.A(_02215_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__inv_2 _18521_ (.A(_02114_),
    .Y(_02219_));
 sky130_fd_sc_hd__o21a_1 _18522_ (.A1(_01922_),
    .A2(_02219_),
    .B1(_02112_),
    .X(_02220_));
 sky130_fd_sc_hd__xnor2_2 _18523_ (.A(_02218_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__a21o_2 _18524_ (.A1(_02138_),
    .A2(_02120_),
    .B1(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__and3_2 _18525_ (.A(_02138_),
    .B(_02120_),
    .C(_02221_),
    .X(_02223_));
 sky130_fd_sc_hd__inv_2 _18526_ (.A(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _18527_ (.A(_02222_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__a21oi_1 _18528_ (.A1(_02125_),
    .A2(_02128_),
    .B1(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__a31o_1 _18529_ (.A1(_02125_),
    .A2(_02128_),
    .A3(_02225_),
    .B1(_05203_),
    .X(_02227_));
 sky130_fd_sc_hd__or2_1 _18530_ (.A(_02226_),
    .B(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__or2_1 _18531_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_02229_));
 sky130_fd_sc_hd__nand2_1 _18532_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_02230_));
 sky130_fd_sc_hd__o21bai_1 _18533_ (.A1(_02132_),
    .A2(_02134_),
    .B1_N(_02133_),
    .Y(_02231_));
 sky130_fd_sc_hd__a21oi_1 _18534_ (.A1(_02229_),
    .A2(_02230_),
    .B1(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__a31o_1 _18535_ (.A1(_02229_),
    .A2(_02230_),
    .A3(_02231_),
    .B1(_05531_),
    .X(_02233_));
 sky130_fd_sc_hd__o21a_1 _18536_ (.A1(_02232_),
    .A2(_02233_),
    .B1(_09817_),
    .X(_02234_));
 sky130_fd_sc_hd__o2bb2a_1 _18537_ (.A1_N(_02228_),
    .A2_N(_02234_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_10036_),
    .X(_00598_));
 sky130_fd_sc_hd__a21bo_1 _18538_ (.A1(_02141_),
    .A2(_02160_),
    .B1_N(_02140_),
    .X(_02235_));
 sky130_fd_sc_hd__o21bai_1 _18539_ (.A1(_02149_),
    .A2(_02156_),
    .B1_N(_02155_),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _18540_ (.A(_01737_),
    .B(_10266_),
    .Y(_02237_));
 sky130_fd_sc_hd__nor2_1 _18541_ (.A(_10238_),
    .B(_09434_),
    .Y(_02238_));
 sky130_fd_sc_hd__xnor2_1 _18542_ (.A(_02237_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _18543_ (.A(_01620_),
    .B(_09292_),
    .Y(_02240_));
 sky130_fd_sc_hd__xnor2_1 _18544_ (.A(_02239_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__o31a_1 _18545_ (.A1(_10248_),
    .A2(_10266_),
    .A3(_02151_),
    .B1(_02045_),
    .X(_02242_));
 sky130_fd_sc_hd__nor2_1 _18546_ (.A(_10248_),
    .B(_01524_),
    .Y(_02243_));
 sky130_fd_sc_hd__xnor2_1 _18547_ (.A(_02151_),
    .B(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__xnor2_1 _18548_ (.A(_02242_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__xor2_1 _18549_ (.A(_02241_),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__xnor2_1 _18550_ (.A(_02144_),
    .B(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__xnor2_1 _18551_ (.A(_02236_),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__xor2_1 _18552_ (.A(_02141_),
    .B(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__xnor2_1 _18553_ (.A(_02235_),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _18554_ (.A(_02193_),
    .B(_02195_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21o_1 _18555_ (.A1(_02184_),
    .A2(_02196_),
    .B1(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__or2b_1 _18556_ (.A(_02159_),
    .B_N(_02143_),
    .X(_02253_));
 sky130_fd_sc_hd__a21bo_1 _18557_ (.A1(_02144_),
    .A2(_02158_),
    .B1_N(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__nor2_1 _18558_ (.A(_10239_),
    .B(_09481_),
    .Y(_02255_));
 sky130_fd_sc_hd__o22a_1 _18559_ (.A1(_10239_),
    .A2(_09350_),
    .B1(_09481_),
    .B2(_10094_),
    .X(_02256_));
 sky130_fd_sc_hd__a21o_1 _18560_ (.A1(_02167_),
    .A2(_02255_),
    .B1(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__nor2_1 _18561_ (.A(_08445_),
    .B(_09704_),
    .Y(_02258_));
 sky130_fd_sc_hd__xnor2_2 _18562_ (.A(_02257_),
    .B(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__or2_1 _18563_ (.A(_08257_),
    .B(_09162_),
    .X(_02260_));
 sky130_fd_sc_hd__or3_1 _18564_ (.A(_01739_),
    .B(_09027_),
    .C(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__o21ai_1 _18565_ (.A1(_01739_),
    .A2(_09027_),
    .B1(_02260_),
    .Y(_02262_));
 sky130_fd_sc_hd__and2_1 _18566_ (.A(_02261_),
    .B(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__nor2_1 _18567_ (.A(_01498_),
    .B(_09215_),
    .Y(_02264_));
 sky130_fd_sc_hd__xnor2_1 _18568_ (.A(_02263_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__a21bo_1 _18569_ (.A1(_02071_),
    .A2(_02172_),
    .B1_N(_02174_),
    .X(_02266_));
 sky130_fd_sc_hd__xnor2_1 _18570_ (.A(_02265_),
    .B(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__xor2_1 _18571_ (.A(_02259_),
    .B(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__a21o_1 _18572_ (.A1(_02039_),
    .A2(_02042_),
    .B1(_02191_),
    .X(_02269_));
 sky130_fd_sc_hd__or2b_1 _18573_ (.A(_02192_),
    .B_N(_02185_),
    .X(_02270_));
 sky130_fd_sc_hd__a21bo_1 _18574_ (.A1(_02188_),
    .A2(_02190_),
    .B1_N(_02187_),
    .X(_02271_));
 sky130_fd_sc_hd__a21bo_1 _18575_ (.A1(_02146_),
    .A2(_02148_),
    .B1_N(_02145_),
    .X(_02272_));
 sky130_fd_sc_hd__nor2_1 _18576_ (.A(_08151_),
    .B(_09138_),
    .Y(_02273_));
 sky130_fd_sc_hd__nor2_1 _18577_ (.A(_09141_),
    .B(_01475_),
    .Y(_02274_));
 sky130_fd_sc_hd__xor2_1 _18578_ (.A(_02273_),
    .B(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_1 _18579_ (.A(_01860_),
    .B(_08423_),
    .Y(_02276_));
 sky130_fd_sc_hd__xor2_1 _18580_ (.A(_02275_),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__and2_1 _18581_ (.A(_02272_),
    .B(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__or2_1 _18582_ (.A(_02272_),
    .B(_02277_),
    .X(_02279_));
 sky130_fd_sc_hd__and2b_1 _18583_ (.A_N(_02278_),
    .B(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__xnor2_1 _18584_ (.A(_02271_),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__a21oi_1 _18585_ (.A1(_02269_),
    .A2(_02270_),
    .B1(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__and3_1 _18586_ (.A(_02269_),
    .B(_02270_),
    .C(_02281_),
    .X(_02283_));
 sky130_fd_sc_hd__nor2_1 _18587_ (.A(_02282_),
    .B(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__xor2_1 _18588_ (.A(_02268_),
    .B(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__xor2_1 _18589_ (.A(_02254_),
    .B(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__xor2_1 _18590_ (.A(_02252_),
    .B(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__xor2_1 _18591_ (.A(_02250_),
    .B(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__nor2_1 _18592_ (.A(_02161_),
    .B(_02162_),
    .Y(_02289_));
 sky130_fd_sc_hd__a21oi_1 _18593_ (.A1(_02163_),
    .A2(_02199_),
    .B1(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__xnor2_1 _18594_ (.A(_02288_),
    .B(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__or2b_1 _18595_ (.A(_02198_),
    .B_N(_02164_),
    .X(_02292_));
 sky130_fd_sc_hd__a21bo_1 _18596_ (.A1(_02166_),
    .A2(_02197_),
    .B1_N(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__or2b_1 _18597_ (.A(_02169_),
    .B_N(_02170_),
    .X(_02294_));
 sky130_fd_sc_hd__a21boi_1 _18598_ (.A1(_02167_),
    .A2(_02168_),
    .B1_N(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__a21oi_1 _18599_ (.A1(_02179_),
    .A2(_02182_),
    .B1(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__and3_1 _18600_ (.A(_02179_),
    .B(_02182_),
    .C(_02295_),
    .X(_02297_));
 sky130_fd_sc_hd__nor2_1 _18601_ (.A(_02296_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__xor2_1 _18602_ (.A(_02293_),
    .B(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__xnor2_1 _18603_ (.A(_02208_),
    .B(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__xor2_1 _18604_ (.A(_02291_),
    .B(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__a21oi_1 _18605_ (.A1(_02204_),
    .A2(_02214_),
    .B1(_02202_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _18606_ (.A(_02301_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__and2_1 _18607_ (.A(_02301_),
    .B(_02302_),
    .X(_02304_));
 sky130_fd_sc_hd__or2_1 _18608_ (.A(_02303_),
    .B(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__a21oi_2 _18609_ (.A1(_02109_),
    .A2(_02213_),
    .B1(_02211_),
    .Y(_02306_));
 sky130_fd_sc_hd__xnor2_2 _18610_ (.A(_02305_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__or2_1 _18611_ (.A(_02215_),
    .B(_02217_),
    .X(_02308_));
 sky130_fd_sc_hd__o21a_1 _18612_ (.A1(_02218_),
    .A2(_02220_),
    .B1(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__nor2_2 _18613_ (.A(_02307_),
    .B(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__and2_1 _18614_ (.A(_02307_),
    .B(_02309_),
    .X(_02311_));
 sky130_fd_sc_hd__or2_2 _18615_ (.A(_02310_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__a311oi_2 _18616_ (.A1(_02125_),
    .A2(_02128_),
    .A3(_02222_),
    .B1(_02223_),
    .C1(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__a31o_1 _18617_ (.A1(_02125_),
    .A2(_02128_),
    .A3(_02222_),
    .B1(_02223_),
    .X(_02314_));
 sky130_fd_sc_hd__a21o_1 _18618_ (.A1(_02312_),
    .A2(_02314_),
    .B1(_05204_),
    .X(_02315_));
 sky130_fd_sc_hd__or2_1 _18619_ (.A(_02313_),
    .B(_02315_),
    .X(_02316_));
 sky130_fd_sc_hd__or2_1 _18620_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_1 _18621_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(_02317_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__a21boi_1 _18623_ (.A1(_02229_),
    .A2(_02231_),
    .B1_N(_02230_),
    .Y(_02320_));
 sky130_fd_sc_hd__xor2_1 _18624_ (.A(_02319_),
    .B(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__a21oi_1 _18625_ (.A1(_09889_),
    .A2(_02321_),
    .B1(_09780_),
    .Y(_02322_));
 sky130_fd_sc_hd__o2bb2a_1 _18626_ (.A1_N(_02316_),
    .A2_N(_02322_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_10036_),
    .X(_00599_));
 sky130_fd_sc_hd__or2b_1 _18627_ (.A(_02291_),
    .B_N(_02300_),
    .X(_02323_));
 sky130_fd_sc_hd__o21a_1 _18628_ (.A1(_02288_),
    .A2(_02290_),
    .B1(_02323_),
    .X(_02324_));
 sky130_fd_sc_hd__xnor2_1 _18629_ (.A(_02296_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21o_1 _18630_ (.A1(_02268_),
    .A2(_02284_),
    .B1(_02282_),
    .X(_02326_));
 sky130_fd_sc_hd__a21oi_1 _18631_ (.A1(_02271_),
    .A2(_02280_),
    .B1(_02278_),
    .Y(_02327_));
 sky130_fd_sc_hd__nor2_1 _18632_ (.A(_08159_),
    .B(_09138_),
    .Y(_02328_));
 sky130_fd_sc_hd__xnor2_1 _18633_ (.A(_02327_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__xnor2_1 _18634_ (.A(_02326_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__a21o_1 _18635_ (.A1(_09429_),
    .A2(_09433_),
    .B1(_08356_),
    .X(_02331_));
 sky130_fd_sc_hd__and2_1 _18636_ (.A(_02273_),
    .B(_02274_),
    .X(_02332_));
 sky130_fd_sc_hd__a21oi_1 _18637_ (.A1(_02275_),
    .A2(_02276_),
    .B1(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__nor2_1 _18638_ (.A(_09141_),
    .B(_08423_),
    .Y(_02334_));
 sky130_fd_sc_hd__xnor2_1 _18639_ (.A(_02333_),
    .B(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__a21o_1 _18640_ (.A1(_09284_),
    .A2(_09287_),
    .B1(_08151_),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_1 _18641_ (.A(_02237_),
    .B(_02238_),
    .Y(_02337_));
 sky130_fd_sc_hd__o31a_1 _18642_ (.A1(_01620_),
    .A2(_09292_),
    .A3(_02239_),
    .B1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _18643_ (.A0(_08418_),
    .A1(_02336_),
    .S(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__xnor2_1 _18644_ (.A(_02335_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__nand2_1 _18645_ (.A(_10094_),
    .B(_09611_),
    .Y(_02341_));
 sky130_fd_sc_hd__xnor2_1 _18646_ (.A(_02340_),
    .B(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__and2_1 _18647_ (.A(_10248_),
    .B(_02150_),
    .X(_02343_));
 sky130_fd_sc_hd__a311o_1 _18648_ (.A1(_02045_),
    .A2(_02150_),
    .A3(_02152_),
    .B1(_02243_),
    .C1(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__a21bo_1 _18649_ (.A1(_02241_),
    .A2(_02245_),
    .B1_N(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__nor2_1 _18650_ (.A(_01739_),
    .B(_09162_),
    .Y(_02346_));
 sky130_fd_sc_hd__xnor2_1 _18651_ (.A(_02345_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__xnor2_1 _18652_ (.A(_02342_),
    .B(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__xnor2_1 _18653_ (.A(_02331_),
    .B(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__xnor2_1 _18654_ (.A(_02330_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__o21a_1 _18655_ (.A1(_02139_),
    .A2(_02248_),
    .B1(_02140_),
    .X(_02351_));
 sky130_fd_sc_hd__and2b_1 _18656_ (.A_N(_02247_),
    .B(_02236_),
    .X(_02352_));
 sky130_fd_sc_hd__a21oi_1 _18657_ (.A1(_02144_),
    .A2(_02246_),
    .B1(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__a21boi_1 _18658_ (.A1(_02263_),
    .A2(_02264_),
    .B1_N(_02261_),
    .Y(_02354_));
 sky130_fd_sc_hd__o22ai_1 _18659_ (.A1(_01860_),
    .A2(_09027_),
    .B1(_09350_),
    .B2(_01498_),
    .Y(_02355_));
 sky130_fd_sc_hd__or4_1 _18660_ (.A(_01498_),
    .B(_01860_),
    .C(_09027_),
    .D(_09350_),
    .X(_02356_));
 sky130_fd_sc_hd__nand2_1 _18661_ (.A(_02355_),
    .B(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__xnor2_1 _18662_ (.A(_02255_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__xnor2_1 _18663_ (.A(_02354_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__nor2_1 _18664_ (.A(_08257_),
    .B(_09215_),
    .Y(_02360_));
 sky130_fd_sc_hd__xnor2_1 _18665_ (.A(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__xnor2_1 _18666_ (.A(_02353_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _18667_ (.A(_02351_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__xnor2_1 _18668_ (.A(_02350_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _18669_ (.A(_02167_),
    .B(_02255_),
    .Y(_02365_));
 sky130_fd_sc_hd__o31a_1 _18670_ (.A1(_08445_),
    .A2(_09704_),
    .A3(_02256_),
    .B1(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__xnor2_1 _18671_ (.A(_02144_),
    .B(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _18672_ (.A(_08047_),
    .B(_09565_),
    .Y(_02368_));
 sky130_fd_sc_hd__or2_1 _18673_ (.A(_01737_),
    .B(_01524_),
    .X(_02369_));
 sky130_fd_sc_hd__and2b_1 _18674_ (.A_N(_02265_),
    .B(_02266_),
    .X(_02370_));
 sky130_fd_sc_hd__a21oi_1 _18675_ (.A1(_02259_),
    .A2(_02267_),
    .B1(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__xnor2_1 _18676_ (.A(_02369_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__xnor2_1 _18677_ (.A(_02368_),
    .B(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__xnor2_1 _18678_ (.A(_02367_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__xnor2_1 _18679_ (.A(_02364_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__and2b_1 _18680_ (.A_N(_02208_),
    .B(_02299_),
    .X(_02376_));
 sky130_fd_sc_hd__a21o_1 _18681_ (.A1(_02293_),
    .A2(_02298_),
    .B1(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__and2b_1 _18682_ (.A_N(_02250_),
    .B(_02287_),
    .X(_02378_));
 sky130_fd_sc_hd__a21oi_1 _18683_ (.A1(_02235_),
    .A2(_02249_),
    .B1(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__xnor2_1 _18684_ (.A(_02377_),
    .B(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__xnor2_1 _18685_ (.A(_02375_),
    .B(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__xnor2_2 _18686_ (.A(_02325_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__o21ba_1 _18687_ (.A1(_02305_),
    .A2(_02306_),
    .B1_N(_02303_),
    .X(_02383_));
 sky130_fd_sc_hd__and2_1 _18688_ (.A(_02254_),
    .B(_02285_),
    .X(_02384_));
 sky130_fd_sc_hd__a21oi_1 _18689_ (.A1(_02252_),
    .A2(_02286_),
    .B1(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__xnor2_2 _18690_ (.A(_02383_),
    .B(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__xor2_4 _18691_ (.A(_02382_),
    .B(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__o21a_1 _18692_ (.A1(_02310_),
    .A2(_02313_),
    .B1(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__or3_1 _18693_ (.A(_02310_),
    .B(_02313_),
    .C(_02387_),
    .X(_02389_));
 sky130_fd_sc_hd__or3b_1 _18694_ (.A(_09889_),
    .B(_02388_),
    .C_N(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__o21ai_1 _18695_ (.A1(_02319_),
    .A2(_02320_),
    .B1(_02318_),
    .Y(_02391_));
 sky130_fd_sc_hd__xor2_1 _18696_ (.A(\rbzero.wall_tracer.trackDistX[11] ),
    .B(\rbzero.wall_tracer.stepDistX[11] ),
    .X(_02392_));
 sky130_fd_sc_hd__xnor2_1 _18697_ (.A(_02391_),
    .B(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__o21a_1 _18698_ (.A1(_05532_),
    .A2(_02393_),
    .B1(_09817_),
    .X(_02394_));
 sky130_fd_sc_hd__o2bb2a_1 _18699_ (.A1_N(_02390_),
    .A2_N(_02394_),
    .B1(\rbzero.wall_tracer.trackDistX[11] ),
    .B2(_10036_),
    .X(_00600_));
 sky130_fd_sc_hd__o21ai_1 _18700_ (.A1(\rbzero.wall_tracer.trackDistY[-12] ),
    .A2(\rbzero.wall_tracer.stepDistY[-12] ),
    .B1(_09807_),
    .Y(_02395_));
 sky130_fd_sc_hd__a21o_1 _18701_ (.A1(\rbzero.wall_tracer.trackDistY[-12] ),
    .A2(\rbzero.wall_tracer.stepDistY[-12] ),
    .B1(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__nand2_1 _18702_ (.A(_09808_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__o21a_2 _18703_ (.A1(_05203_),
    .A2(_09283_),
    .B1(_05282_),
    .X(_02398_));
 sky130_fd_sc_hd__buf_4 _18704_ (.A(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _18705_ (.A0(\rbzero.wall_tracer.trackDistY[-12] ),
    .A1(_02397_),
    .S(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__clkbuf_1 _18706_ (.A(_02400_),
    .X(_00601_));
 sky130_fd_sc_hd__or2_1 _18707_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_02401_));
 sky130_fd_sc_hd__nand2_1 _18708_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_02402_));
 sky130_fd_sc_hd__and4_1 _18709_ (.A(\rbzero.wall_tracer.trackDistY[-12] ),
    .B(\rbzero.wall_tracer.stepDistY[-12] ),
    .C(_02401_),
    .D(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__a22oi_1 _18710_ (.A1(\rbzero.wall_tracer.trackDistY[-12] ),
    .A2(\rbzero.wall_tracer.stepDistY[-12] ),
    .B1(_02401_),
    .B2(_02402_),
    .Y(_02404_));
 sky130_fd_sc_hd__o31a_1 _18711_ (.A1(_05532_),
    .A2(_02403_),
    .A3(_02404_),
    .B1(_02399_),
    .X(_02405_));
 sky130_fd_sc_hd__buf_4 _18712_ (.A(_02398_),
    .X(_02406_));
 sky130_fd_sc_hd__o2bb2a_1 _18713_ (.A1_N(_02405_),
    .A2_N(_09819_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .B2(_02406_),
    .X(_00602_));
 sky130_fd_sc_hd__a21oi_1 _18714_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(\rbzero.wall_tracer.stepDistY[-11] ),
    .B1(_02403_),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_1 _18715_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_02408_));
 sky130_fd_sc_hd__and2_1 _18716_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_02409_));
 sky130_fd_sc_hd__nor3_1 _18717_ (.A(_02407_),
    .B(_02408_),
    .C(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__o21a_1 _18718_ (.A1(_02408_),
    .A2(_02409_),
    .B1(_02407_),
    .X(_02411_));
 sky130_fd_sc_hd__o31ai_1 _18719_ (.A1(_09863_),
    .A2(_02410_),
    .A3(_02411_),
    .B1(_09827_),
    .Y(_02412_));
 sky130_fd_sc_hd__mux2_1 _18720_ (.A0(\rbzero.wall_tracer.trackDistY[-10] ),
    .A1(_02412_),
    .S(_02399_),
    .X(_02413_));
 sky130_fd_sc_hd__clkbuf_1 _18721_ (.A(_02413_),
    .X(_00603_));
 sky130_fd_sc_hd__or2_1 _18722_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_02414_));
 sky130_fd_sc_hd__nand2_1 _18723_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_02415_));
 sky130_fd_sc_hd__o21bai_1 _18724_ (.A1(_02407_),
    .A2(_02408_),
    .B1_N(_02409_),
    .Y(_02416_));
 sky130_fd_sc_hd__and3_1 _18725_ (.A(_02414_),
    .B(_02415_),
    .C(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__a21oi_1 _18726_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_02416_),
    .Y(_02418_));
 sky130_fd_sc_hd__o31ai_1 _18727_ (.A1(_09863_),
    .A2(_02417_),
    .A3(_02418_),
    .B1(_09835_),
    .Y(_02419_));
 sky130_fd_sc_hd__mux2_1 _18728_ (.A0(\rbzero.wall_tracer.trackDistY[-9] ),
    .A1(_02419_),
    .S(_02399_),
    .X(_02420_));
 sky130_fd_sc_hd__clkbuf_1 _18729_ (.A(_02420_),
    .X(_00604_));
 sky130_fd_sc_hd__nor2_1 _18730_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_02421_));
 sky130_fd_sc_hd__and2_1 _18731_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_02422_));
 sky130_fd_sc_hd__a21boi_1 _18732_ (.A1(_02414_),
    .A2(_02416_),
    .B1_N(_02415_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor3_1 _18733_ (.A(_02421_),
    .B(_02422_),
    .C(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__o21a_1 _18734_ (.A1(_02421_),
    .A2(_02422_),
    .B1(_02423_),
    .X(_02425_));
 sky130_fd_sc_hd__o31ai_1 _18735_ (.A1(_09863_),
    .A2(_02424_),
    .A3(_02425_),
    .B1(_09843_),
    .Y(_02426_));
 sky130_fd_sc_hd__mux2_1 _18736_ (.A0(\rbzero.wall_tracer.trackDistY[-8] ),
    .A1(_02426_),
    .S(_02399_),
    .X(_02427_));
 sky130_fd_sc_hd__clkbuf_1 _18737_ (.A(_02427_),
    .X(_00605_));
 sky130_fd_sc_hd__or2_1 _18738_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .X(_02428_));
 sky130_fd_sc_hd__nand2_1 _18739_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02429_));
 sky130_fd_sc_hd__o21bai_1 _18740_ (.A1(_02421_),
    .A2(_02423_),
    .B1_N(_02422_),
    .Y(_02430_));
 sky130_fd_sc_hd__a21oi_1 _18741_ (.A1(_02428_),
    .A2(_02429_),
    .B1(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__a31o_1 _18742_ (.A1(_02428_),
    .A2(_02429_),
    .A3(_02430_),
    .B1(_05531_),
    .X(_02432_));
 sky130_fd_sc_hd__o21ai_1 _18743_ (.A1(_02431_),
    .A2(_02432_),
    .B1(_09851_),
    .Y(_02433_));
 sky130_fd_sc_hd__mux2_1 _18744_ (.A0(\rbzero.wall_tracer.trackDistY[-7] ),
    .A1(_02433_),
    .S(_02399_),
    .X(_02434_));
 sky130_fd_sc_hd__clkbuf_1 _18745_ (.A(_02434_),
    .X(_00606_));
 sky130_fd_sc_hd__nor2_1 _18746_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_02435_));
 sky130_fd_sc_hd__and2_1 _18747_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_02436_));
 sky130_fd_sc_hd__a21boi_1 _18748_ (.A1(_02428_),
    .A2(_02430_),
    .B1_N(_02429_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor3_1 _18749_ (.A(_02435_),
    .B(_02436_),
    .C(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__o21a_1 _18750_ (.A1(_02435_),
    .A2(_02436_),
    .B1(_02437_),
    .X(_02439_));
 sky130_fd_sc_hd__o31ai_1 _18751_ (.A1(_09863_),
    .A2(_02438_),
    .A3(_02439_),
    .B1(_09860_),
    .Y(_02440_));
 sky130_fd_sc_hd__buf_6 _18752_ (.A(_02398_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _18753_ (.A0(\rbzero.wall_tracer.trackDistY[-6] ),
    .A1(_02440_),
    .S(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__clkbuf_1 _18754_ (.A(_02442_),
    .X(_00607_));
 sky130_fd_sc_hd__or2_1 _18755_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .X(_02443_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02444_));
 sky130_fd_sc_hd__o21bai_1 _18757_ (.A1(_02435_),
    .A2(_02437_),
    .B1_N(_02436_),
    .Y(_02445_));
 sky130_fd_sc_hd__and3_1 _18758_ (.A(_02443_),
    .B(_02444_),
    .C(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__a21oi_1 _18759_ (.A1(_02443_),
    .A2(_02444_),
    .B1(_02445_),
    .Y(_02447_));
 sky130_fd_sc_hd__o31ai_1 _18760_ (.A1(_09863_),
    .A2(_02446_),
    .A3(_02447_),
    .B1(_09869_),
    .Y(_02448_));
 sky130_fd_sc_hd__mux2_1 _18761_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(_02448_),
    .S(_02441_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_1 _18762_ (.A(_02449_),
    .X(_00608_));
 sky130_fd_sc_hd__nor2_1 _18763_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02450_));
 sky130_fd_sc_hd__nand2_1 _18764_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02451_));
 sky130_fd_sc_hd__or2b_1 _18765_ (.A(_02450_),
    .B_N(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__a21boi_1 _18766_ (.A1(_02443_),
    .A2(_02445_),
    .B1_N(_02444_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_1 _18767_ (.A(_02452_),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__o21ai_1 _18768_ (.A1(_09812_),
    .A2(_02454_),
    .B1(_09877_),
    .Y(_02455_));
 sky130_fd_sc_hd__mux2_1 _18769_ (.A0(\rbzero.wall_tracer.trackDistY[-4] ),
    .A1(_02455_),
    .S(_02441_),
    .X(_02456_));
 sky130_fd_sc_hd__clkbuf_1 _18770_ (.A(_02456_),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _18771_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_1 _18772_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02458_));
 sky130_fd_sc_hd__o21ai_1 _18773_ (.A1(_02450_),
    .A2(_02453_),
    .B1(_02451_),
    .Y(_02459_));
 sky130_fd_sc_hd__and3_1 _18774_ (.A(_02457_),
    .B(_02458_),
    .C(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__a21oi_1 _18775_ (.A1(_02457_),
    .A2(_02458_),
    .B1(_02459_),
    .Y(_02461_));
 sky130_fd_sc_hd__o31ai_1 _18776_ (.A1(_09863_),
    .A2(_02460_),
    .A3(_02461_),
    .B1(_09885_),
    .Y(_02462_));
 sky130_fd_sc_hd__mux2_1 _18777_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(_02462_),
    .S(_02441_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _18778_ (.A(_02463_),
    .X(_00610_));
 sky130_fd_sc_hd__nand2_1 _18779_ (.A(_09812_),
    .B(_09597_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_1 _18780_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02465_));
 sky130_fd_sc_hd__and2_1 _18781_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_02466_));
 sky130_fd_sc_hd__a21boi_1 _18782_ (.A1(_02457_),
    .A2(_02459_),
    .B1_N(_02458_),
    .Y(_02467_));
 sky130_fd_sc_hd__o21a_1 _18783_ (.A1(_02465_),
    .A2(_02466_),
    .B1(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__or3_1 _18784_ (.A(_02465_),
    .B(_02466_),
    .C(_02467_),
    .X(_02469_));
 sky130_fd_sc_hd__or3b_1 _18785_ (.A(_02468_),
    .B(_05531_),
    .C_N(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__and3_1 _18786_ (.A(_02464_),
    .B(_02398_),
    .C(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__o21ba_1 _18787_ (.A1(\rbzero.wall_tracer.trackDistY[-2] ),
    .A2(_02406_),
    .B1_N(_02471_),
    .X(_00611_));
 sky130_fd_sc_hd__nor2_1 _18788_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02472_));
 sky130_fd_sc_hd__and2_1 _18789_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(_02473_));
 sky130_fd_sc_hd__nand2_1 _18790_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02474_));
 sky130_fd_sc_hd__o211ai_1 _18791_ (.A1(_02472_),
    .A2(_02473_),
    .B1(_02474_),
    .C1(_02469_),
    .Y(_02475_));
 sky130_fd_sc_hd__a211o_1 _18792_ (.A1(_02474_),
    .A2(_02469_),
    .B1(_02472_),
    .C1(_02473_),
    .X(_02476_));
 sky130_fd_sc_hd__a31o_1 _18793_ (.A1(_05204_),
    .A2(_02475_),
    .A3(_02476_),
    .B1(_09897_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _18794_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(_02477_),
    .S(_02441_),
    .X(_02478_));
 sky130_fd_sc_hd__clkbuf_1 _18795_ (.A(_02478_),
    .X(_00612_));
 sky130_fd_sc_hd__nand2_1 _18796_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _18797_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_02480_));
 sky130_fd_sc_hd__nor2_1 _18798_ (.A(_05257_),
    .B(_08200_),
    .Y(_02481_));
 sky130_fd_sc_hd__a211o_1 _18799_ (.A1(_02479_),
    .A2(_02476_),
    .B1(_02480_),
    .C1(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__inv_2 _18800_ (.A(_02482_),
    .Y(_02483_));
 sky130_fd_sc_hd__o211a_1 _18801_ (.A1(_02480_),
    .A2(_02481_),
    .B1(_02479_),
    .C1(_02476_),
    .X(_02484_));
 sky130_fd_sc_hd__o31a_1 _18802_ (.A1(_05532_),
    .A2(_02483_),
    .A3(_02484_),
    .B1(_02399_),
    .X(_02485_));
 sky130_fd_sc_hd__o2bb2a_1 _18803_ (.A1_N(_02485_),
    .A2_N(_10028_),
    .B1(\rbzero.wall_tracer.trackDistY[0] ),
    .B2(_02406_),
    .X(_00613_));
 sky130_fd_sc_hd__or2_1 _18804_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_02486_));
 sky130_fd_sc_hd__nand2_1 _18805_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_02487_));
 sky130_fd_sc_hd__a211o_1 _18806_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_02481_),
    .C1(_02483_),
    .X(_02488_));
 sky130_fd_sc_hd__o211ai_2 _18807_ (.A1(_02481_),
    .A2(_02483_),
    .B1(_02486_),
    .C1(_02487_),
    .Y(_02489_));
 sky130_fd_sc_hd__a31o_1 _18808_ (.A1(_05204_),
    .A2(_02488_),
    .A3(_02489_),
    .B1(_10173_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _18809_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(_02490_),
    .S(_02441_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _18810_ (.A(_02491_),
    .X(_00614_));
 sky130_fd_sc_hd__nor2_1 _18811_ (.A(_05254_),
    .B(_08186_),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2_1 _18812_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_02493_));
 sky130_fd_sc_hd__a211oi_1 _18813_ (.A1(_02487_),
    .A2(_02489_),
    .B1(_02492_),
    .C1(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__o211a_1 _18814_ (.A1(_02492_),
    .A2(_02493_),
    .B1(_02487_),
    .C1(_02489_),
    .X(_02495_));
 sky130_fd_sc_hd__o31a_1 _18815_ (.A1(_05532_),
    .A2(_02494_),
    .A3(_02495_),
    .B1(_02399_),
    .X(_02496_));
 sky130_fd_sc_hd__o2bb2a_1 _18816_ (.A1_N(_02496_),
    .A2_N(_01438_),
    .B1(\rbzero.wall_tracer.trackDistY[2] ),
    .B2(_02406_),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_1 _18817_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_02497_));
 sky130_fd_sc_hd__or2_1 _18818_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_02498_));
 sky130_fd_sc_hd__nand2_1 _18819_ (.A(_02497_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__or2_1 _18820_ (.A(_02492_),
    .B(_02494_),
    .X(_02500_));
 sky130_fd_sc_hd__xnor2_1 _18821_ (.A(_02499_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__a21boi_1 _18822_ (.A1(_09889_),
    .A2(_02501_),
    .B1_N(_02399_),
    .Y(_02502_));
 sky130_fd_sc_hd__o2bb2a_1 _18823_ (.A1_N(_02502_),
    .A2_N(_01553_),
    .B1(\rbzero.wall_tracer.trackDistY[3] ),
    .B2(_02406_),
    .X(_00616_));
 sky130_fd_sc_hd__nor2_1 _18824_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_02503_));
 sky130_fd_sc_hd__and2_1 _18825_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_02504_));
 sky130_fd_sc_hd__a21boi_1 _18826_ (.A1(_02498_),
    .A2(_02500_),
    .B1_N(_02497_),
    .Y(_02505_));
 sky130_fd_sc_hd__nor3_1 _18827_ (.A(_02503_),
    .B(_02504_),
    .C(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__o21a_1 _18828_ (.A1(_02503_),
    .A2(_02504_),
    .B1(_02505_),
    .X(_02507_));
 sky130_fd_sc_hd__o31ai_1 _18829_ (.A1(_09863_),
    .A2(_02506_),
    .A3(_02507_),
    .B1(_01677_),
    .Y(_02508_));
 sky130_fd_sc_hd__mux2_1 _18830_ (.A0(\rbzero.wall_tracer.trackDistY[4] ),
    .A1(_02508_),
    .S(_02441_),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_1 _18831_ (.A(_02509_),
    .X(_00617_));
 sky130_fd_sc_hd__or2_1 _18832_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_02510_));
 sky130_fd_sc_hd__nand2_1 _18833_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_02511_));
 sky130_fd_sc_hd__o21bai_1 _18834_ (.A1(_02503_),
    .A2(_02505_),
    .B1_N(_02504_),
    .Y(_02512_));
 sky130_fd_sc_hd__a21oi_1 _18835_ (.A1(_02510_),
    .A2(_02511_),
    .B1(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__a31o_1 _18836_ (.A1(_02510_),
    .A2(_02511_),
    .A3(_02512_),
    .B1(_04016_),
    .X(_02514_));
 sky130_fd_sc_hd__o21ai_1 _18837_ (.A1(_02513_),
    .A2(_02514_),
    .B1(_01792_),
    .Y(_02515_));
 sky130_fd_sc_hd__mux2_1 _18838_ (.A0(\rbzero.wall_tracer.trackDistY[5] ),
    .A1(_02515_),
    .S(_02441_),
    .X(_02516_));
 sky130_fd_sc_hd__clkbuf_1 _18839_ (.A(_02516_),
    .X(_00618_));
 sky130_fd_sc_hd__nor2_1 _18840_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02517_));
 sky130_fd_sc_hd__and2_1 _18841_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .X(_02518_));
 sky130_fd_sc_hd__a21boi_1 _18842_ (.A1(_02510_),
    .A2(_02512_),
    .B1_N(_02511_),
    .Y(_02519_));
 sky130_fd_sc_hd__o21ai_1 _18843_ (.A1(_02517_),
    .A2(_02518_),
    .B1(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__o31a_1 _18844_ (.A1(_02517_),
    .A2(_02518_),
    .A3(_02519_),
    .B1(_09807_),
    .X(_02521_));
 sky130_fd_sc_hd__a21bo_1 _18845_ (.A1(_02520_),
    .A2(_02521_),
    .B1_N(_01908_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _18846_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(_02522_),
    .S(_02441_),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _18847_ (.A(_02523_),
    .X(_00619_));
 sky130_fd_sc_hd__or2_1 _18848_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .X(_02524_));
 sky130_fd_sc_hd__nand2_1 _18849_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02525_));
 sky130_fd_sc_hd__o21bai_1 _18850_ (.A1(_02517_),
    .A2(_02519_),
    .B1_N(_02518_),
    .Y(_02526_));
 sky130_fd_sc_hd__a21oi_1 _18851_ (.A1(_02524_),
    .A2(_02525_),
    .B1(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__a31o_1 _18852_ (.A1(_02524_),
    .A2(_02525_),
    .A3(_02526_),
    .B1(_05531_),
    .X(_02528_));
 sky130_fd_sc_hd__o21a_1 _18853_ (.A1(_02527_),
    .A2(_02528_),
    .B1(_02406_),
    .X(_02529_));
 sky130_fd_sc_hd__o2bb2a_1 _18854_ (.A1_N(_02529_),
    .A2_N(_02016_),
    .B1(\rbzero.wall_tracer.trackDistY[7] ),
    .B2(_02406_),
    .X(_00620_));
 sky130_fd_sc_hd__nor2_1 _18855_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02530_));
 sky130_fd_sc_hd__and2_1 _18856_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_02531_));
 sky130_fd_sc_hd__a21boi_1 _18857_ (.A1(_02524_),
    .A2(_02526_),
    .B1_N(_02525_),
    .Y(_02532_));
 sky130_fd_sc_hd__o21ai_1 _18858_ (.A1(_02530_),
    .A2(_02531_),
    .B1(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__o31a_1 _18859_ (.A1(_02530_),
    .A2(_02531_),
    .A3(_02532_),
    .B1(_05203_),
    .X(_02534_));
 sky130_fd_sc_hd__a22o_1 _18860_ (.A1(_02128_),
    .A2(_02130_),
    .B1(_02533_),
    .B2(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _18861_ (.A0(\rbzero.wall_tracer.trackDistY[8] ),
    .A1(_02535_),
    .S(_02441_),
    .X(_02536_));
 sky130_fd_sc_hd__clkbuf_1 _18862_ (.A(_02536_),
    .X(_00621_));
 sky130_fd_sc_hd__or2_1 _18863_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_02537_));
 sky130_fd_sc_hd__nand2_1 _18864_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_02538_));
 sky130_fd_sc_hd__o21bai_1 _18865_ (.A1(_02530_),
    .A2(_02532_),
    .B1_N(_02531_),
    .Y(_02539_));
 sky130_fd_sc_hd__a21oi_1 _18866_ (.A1(_02537_),
    .A2(_02538_),
    .B1(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__a31o_1 _18867_ (.A1(_02537_),
    .A2(_02538_),
    .A3(_02539_),
    .B1(_04016_),
    .X(_02541_));
 sky130_fd_sc_hd__o21ai_1 _18868_ (.A1(_02540_),
    .A2(_02541_),
    .B1(_02228_),
    .Y(_02542_));
 sky130_fd_sc_hd__mux2_1 _18869_ (.A0(\rbzero.wall_tracer.trackDistY[9] ),
    .A1(_02542_),
    .S(_02398_),
    .X(_02543_));
 sky130_fd_sc_hd__clkbuf_1 _18870_ (.A(_02543_),
    .X(_00622_));
 sky130_fd_sc_hd__or2_1 _18871_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .X(_02544_));
 sky130_fd_sc_hd__nand2_1 _18872_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2_1 _18873_ (.A(_02544_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__a21boi_1 _18874_ (.A1(_02537_),
    .A2(_02539_),
    .B1_N(_02538_),
    .Y(_02547_));
 sky130_fd_sc_hd__xnor2_1 _18875_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21a_1 _18876_ (.A1(_05532_),
    .A2(_02548_),
    .B1(_02406_),
    .X(_02549_));
 sky130_fd_sc_hd__o2bb2a_1 _18877_ (.A1_N(_02549_),
    .A2_N(_02316_),
    .B1(\rbzero.wall_tracer.trackDistY[10] ),
    .B2(_02406_),
    .X(_00623_));
 sky130_fd_sc_hd__o21ai_1 _18878_ (.A1(_02546_),
    .A2(_02547_),
    .B1(_02545_),
    .Y(_02550_));
 sky130_fd_sc_hd__xor2_1 _18879_ (.A(\rbzero.wall_tracer.trackDistY[11] ),
    .B(\rbzero.wall_tracer.stepDistY[11] ),
    .X(_02551_));
 sky130_fd_sc_hd__xnor2_1 _18880_ (.A(_02550_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__o21a_1 _18881_ (.A1(_05532_),
    .A2(_02552_),
    .B1(_02399_),
    .X(_02553_));
 sky130_fd_sc_hd__o2bb2a_1 _18882_ (.A1_N(_02553_),
    .A2_N(_02390_),
    .B1(\rbzero.wall_tracer.trackDistY[11] ),
    .B2(_02406_),
    .X(_00624_));
 sky130_fd_sc_hd__and4bb_1 _18883_ (.A_N(\rbzero.spi_registers.spi_cmd[1] ),
    .B_N(\rbzero.spi_registers.spi_cmd[3] ),
    .C(\rbzero.spi_registers.spi_cmd[2] ),
    .D(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02554_));
 sky130_fd_sc_hd__and3_1 _18884_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_03480_),
    .C(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _18885_ (.A0(\rbzero.spi_registers.new_vinf ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__clkbuf_1 _18886_ (.A(_02556_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_2 _18887_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_03555_),
    .Y(_02557_));
 sky130_fd_sc_hd__nor2b_2 _18888_ (.A(\rbzero.spi_registers.sclk_buffer[2] ),
    .B_N(\rbzero.spi_registers.sclk_buffer[1] ),
    .Y(_02558_));
 sky130_fd_sc_hd__inv_2 _18889_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _18890_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .Y(_02560_));
 sky130_fd_sc_hd__or2_1 _18891_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02561_));
 sky130_fd_sc_hd__or3b_1 _18892_ (.A(_02561_),
    .B(\rbzero.spi_registers.spi_cmd[3] ),
    .C_N(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_02562_));
 sky130_fd_sc_hd__inv_2 _18893_ (.A(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _18894_ (.A(_02560_),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__a21o_1 _18895_ (.A1(\rbzero.spi_registers.spi_cmd[1] ),
    .A2(\rbzero.spi_registers.spi_cmd[0] ),
    .B1(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__xnor2_1 _18896_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__or3_1 _18897_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .C(\rbzero.spi_registers.spi_counter[4] ),
    .X(_02567_));
 sky130_fd_sc_hd__a21oi_1 _18898_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02564_),
    .B1(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__and3_1 _18899_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .C(_02560_),
    .X(_02569_));
 sky130_fd_sc_hd__xnor2_1 _18900_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__o21a_1 _18901_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(_02564_),
    .B1(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__o2111a_1 _18902_ (.A1(_02559_),
    .A2(\rbzero.spi_registers.spi_counter[0] ),
    .B1(_02566_),
    .C1(_02568_),
    .D1(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__nand2_1 _18903_ (.A(_02558_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__and2_1 _18904_ (.A(_02557_),
    .B(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__or2_1 _18905_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .B(_02558_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_1 _18906_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .B(_02558_),
    .Y(_02576_));
 sky130_fd_sc_hd__and3_1 _18907_ (.A(_02574_),
    .B(_02575_),
    .C(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__clkbuf_1 _18908_ (.A(_02577_),
    .X(_00626_));
 sky130_fd_sc_hd__xnor2_1 _18909_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(_02576_),
    .Y(_02578_));
 sky130_fd_sc_hd__and3_1 _18910_ (.A(_02557_),
    .B(_02573_),
    .C(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__clkbuf_1 _18911_ (.A(_02579_),
    .X(_00627_));
 sky130_fd_sc_hd__and4_1 _18912_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_counter[1] ),
    .C(\rbzero.spi_registers.spi_counter[0] ),
    .D(_02558_),
    .X(_02580_));
 sky130_fd_sc_hd__a31o_1 _18913_ (.A1(\rbzero.spi_registers.spi_counter[1] ),
    .A2(\rbzero.spi_registers.spi_counter[0] ),
    .A3(_02558_),
    .B1(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02581_));
 sky130_fd_sc_hd__and3b_1 _18914_ (.A_N(_02580_),
    .B(_02581_),
    .C(_02574_),
    .X(_02582_));
 sky130_fd_sc_hd__clkbuf_1 _18915_ (.A(_02582_),
    .X(_00628_));
 sky130_fd_sc_hd__and2_1 _18916_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02580_),
    .X(_02583_));
 sky130_fd_sc_hd__or2_1 _18917_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02580_),
    .X(_02584_));
 sky130_fd_sc_hd__and3b_1 _18918_ (.A_N(_02583_),
    .B(_02584_),
    .C(_02574_),
    .X(_02585_));
 sky130_fd_sc_hd__clkbuf_1 _18919_ (.A(_02585_),
    .X(_00629_));
 sky130_fd_sc_hd__nand2_1 _18920_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02583_),
    .Y(_02586_));
 sky130_fd_sc_hd__or2_1 _18921_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02583_),
    .X(_02587_));
 sky130_fd_sc_hd__and3_1 _18922_ (.A(_02574_),
    .B(_02586_),
    .C(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__clkbuf_1 _18923_ (.A(_02588_),
    .X(_00630_));
 sky130_fd_sc_hd__and3_1 _18924_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(\rbzero.spi_registers.spi_counter[4] ),
    .C(_02583_),
    .X(_02589_));
 sky130_fd_sc_hd__a31o_1 _18925_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(\rbzero.spi_registers.spi_counter[3] ),
    .A3(_02580_),
    .B1(\rbzero.spi_registers.spi_counter[5] ),
    .X(_02590_));
 sky130_fd_sc_hd__and3b_1 _18926_ (.A_N(_02589_),
    .B(_02557_),
    .C(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__clkbuf_1 _18927_ (.A(_02591_),
    .X(_00631_));
 sky130_fd_sc_hd__o21ai_1 _18928_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02589_),
    .B1(_02557_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _18929_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02589_),
    .B1(_02592_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _18930_ (.A(\rbzero.pov.spi_done ),
    .B(_03480_),
    .Y(_02593_));
 sky130_fd_sc_hd__buf_4 _18931_ (.A(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__clkbuf_4 _18932_ (.A(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _18933_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.ready_buffer[0] ),
    .S(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__clkbuf_1 _18934_ (.A(_02596_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _18935_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.ready_buffer[1] ),
    .S(_02595_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_1 _18936_ (.A(_02597_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _18937_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.ready_buffer[2] ),
    .S(_02595_),
    .X(_02598_));
 sky130_fd_sc_hd__clkbuf_1 _18938_ (.A(_02598_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _18939_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.ready_buffer[3] ),
    .S(_02595_),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_1 _18940_ (.A(_02599_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _18941_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.ready_buffer[4] ),
    .S(_02595_),
    .X(_02600_));
 sky130_fd_sc_hd__clkbuf_1 _18942_ (.A(_02600_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _18943_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.ready_buffer[5] ),
    .S(_02595_),
    .X(_02601_));
 sky130_fd_sc_hd__clkbuf_1 _18944_ (.A(_02601_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _18945_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.ready_buffer[6] ),
    .S(_02595_),
    .X(_02602_));
 sky130_fd_sc_hd__clkbuf_1 _18946_ (.A(_02602_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _18947_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.ready_buffer[7] ),
    .S(_02595_),
    .X(_02603_));
 sky130_fd_sc_hd__clkbuf_1 _18948_ (.A(_02603_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _18949_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.ready_buffer[8] ),
    .S(_02595_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_1 _18950_ (.A(_02604_),
    .X(_00641_));
 sky130_fd_sc_hd__clkbuf_4 _18951_ (.A(_02594_),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _18952_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.ready_buffer[9] ),
    .S(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__clkbuf_1 _18953_ (.A(_02606_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _18954_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.ready_buffer[10] ),
    .S(_02605_),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_1 _18955_ (.A(_02607_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _18956_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.ready_buffer[11] ),
    .S(_02605_),
    .X(_02608_));
 sky130_fd_sc_hd__clkbuf_1 _18957_ (.A(_02608_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _18958_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.ready_buffer[12] ),
    .S(_02605_),
    .X(_02609_));
 sky130_fd_sc_hd__clkbuf_1 _18959_ (.A(_02609_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _18960_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.ready_buffer[13] ),
    .S(_02605_),
    .X(_02610_));
 sky130_fd_sc_hd__clkbuf_1 _18961_ (.A(_02610_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _18962_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.ready_buffer[14] ),
    .S(_02605_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_1 _18963_ (.A(_02611_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18964_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.ready_buffer[15] ),
    .S(_02605_),
    .X(_02612_));
 sky130_fd_sc_hd__clkbuf_1 _18965_ (.A(_02612_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _18966_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.ready_buffer[16] ),
    .S(_02605_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_1 _18967_ (.A(_02613_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18968_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.ready_buffer[17] ),
    .S(_02605_),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_1 _18969_ (.A(_02614_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18970_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.ready_buffer[18] ),
    .S(_02605_),
    .X(_02615_));
 sky130_fd_sc_hd__clkbuf_1 _18971_ (.A(_02615_),
    .X(_00651_));
 sky130_fd_sc_hd__clkbuf_4 _18972_ (.A(_02594_),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _18973_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.ready_buffer[19] ),
    .S(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__clkbuf_1 _18974_ (.A(_02617_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18975_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.ready_buffer[20] ),
    .S(_02616_),
    .X(_02618_));
 sky130_fd_sc_hd__clkbuf_1 _18976_ (.A(_02618_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18977_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.ready_buffer[21] ),
    .S(_02616_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _18978_ (.A(_02619_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18979_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.ready_buffer[22] ),
    .S(_02616_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_1 _18980_ (.A(_02620_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _18981_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.ready_buffer[23] ),
    .S(_02616_),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_1 _18982_ (.A(_02621_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18983_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.ready_buffer[24] ),
    .S(_02616_),
    .X(_02622_));
 sky130_fd_sc_hd__clkbuf_1 _18984_ (.A(_02622_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _18985_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.ready_buffer[25] ),
    .S(_02616_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _18986_ (.A(_02623_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _18987_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.ready_buffer[26] ),
    .S(_02616_),
    .X(_02624_));
 sky130_fd_sc_hd__clkbuf_1 _18988_ (.A(_02624_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18989_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.ready_buffer[27] ),
    .S(_02616_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _18990_ (.A(_02625_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18991_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.ready_buffer[28] ),
    .S(_02616_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _18992_ (.A(_02626_),
    .X(_00661_));
 sky130_fd_sc_hd__buf_4 _18993_ (.A(_02594_),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _18994_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.ready_buffer[29] ),
    .S(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_1 _18995_ (.A(_02628_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _18996_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.ready_buffer[30] ),
    .S(_02627_),
    .X(_02629_));
 sky130_fd_sc_hd__clkbuf_1 _18997_ (.A(_02629_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _18998_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.ready_buffer[31] ),
    .S(_02627_),
    .X(_02630_));
 sky130_fd_sc_hd__clkbuf_1 _18999_ (.A(_02630_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _19000_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.ready_buffer[32] ),
    .S(_02627_),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_1 _19001_ (.A(_02631_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _19002_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.ready_buffer[33] ),
    .S(_02627_),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_1 _19003_ (.A(_02632_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _19004_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.ready_buffer[34] ),
    .S(_02627_),
    .X(_02633_));
 sky130_fd_sc_hd__clkbuf_1 _19005_ (.A(_02633_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _19006_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.ready_buffer[35] ),
    .S(_02627_),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _19007_ (.A(_02634_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _19008_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.ready_buffer[36] ),
    .S(_02627_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _19009_ (.A(_02635_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _19010_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.ready_buffer[37] ),
    .S(_02627_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_1 _19011_ (.A(_02636_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _19012_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.ready_buffer[38] ),
    .S(_02627_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_1 _19013_ (.A(_02637_),
    .X(_00671_));
 sky130_fd_sc_hd__buf_4 _19014_ (.A(_02594_),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _19015_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.ready_buffer[39] ),
    .S(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__clkbuf_1 _19016_ (.A(_02639_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _19017_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.ready_buffer[40] ),
    .S(_02638_),
    .X(_02640_));
 sky130_fd_sc_hd__clkbuf_1 _19018_ (.A(_02640_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _19019_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.ready_buffer[41] ),
    .S(_02638_),
    .X(_02641_));
 sky130_fd_sc_hd__clkbuf_1 _19020_ (.A(_02641_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _19021_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.ready_buffer[42] ),
    .S(_02638_),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_1 _19022_ (.A(_02642_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _19023_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.ready_buffer[43] ),
    .S(_02638_),
    .X(_02643_));
 sky130_fd_sc_hd__clkbuf_1 _19024_ (.A(_02643_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _19025_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_02638_),
    .X(_02644_));
 sky130_fd_sc_hd__clkbuf_1 _19026_ (.A(_02644_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _19027_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.ready_buffer[45] ),
    .S(_02638_),
    .X(_02645_));
 sky130_fd_sc_hd__clkbuf_1 _19028_ (.A(_02645_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _19029_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.ready_buffer[46] ),
    .S(_02638_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_1 _19030_ (.A(_02646_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _19031_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.ready_buffer[47] ),
    .S(_02638_),
    .X(_02647_));
 sky130_fd_sc_hd__clkbuf_1 _19032_ (.A(_02647_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _19033_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.ready_buffer[48] ),
    .S(_02638_),
    .X(_02648_));
 sky130_fd_sc_hd__clkbuf_1 _19034_ (.A(_02648_),
    .X(_00681_));
 sky130_fd_sc_hd__clkbuf_4 _19035_ (.A(_02593_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _19036_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.ready_buffer[49] ),
    .S(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__clkbuf_1 _19037_ (.A(_02650_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _19038_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.ready_buffer[50] ),
    .S(_02649_),
    .X(_02651_));
 sky130_fd_sc_hd__clkbuf_1 _19039_ (.A(_02651_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _19040_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.ready_buffer[51] ),
    .S(_02649_),
    .X(_02652_));
 sky130_fd_sc_hd__clkbuf_1 _19041_ (.A(_02652_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _19042_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.ready_buffer[52] ),
    .S(_02649_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_1 _19043_ (.A(_02653_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _19044_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.ready_buffer[53] ),
    .S(_02649_),
    .X(_02654_));
 sky130_fd_sc_hd__clkbuf_1 _19045_ (.A(_02654_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _19046_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.ready_buffer[54] ),
    .S(_02649_),
    .X(_02655_));
 sky130_fd_sc_hd__clkbuf_1 _19047_ (.A(_02655_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _19048_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.ready_buffer[55] ),
    .S(_02649_),
    .X(_02656_));
 sky130_fd_sc_hd__clkbuf_1 _19049_ (.A(_02656_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _19050_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.ready_buffer[56] ),
    .S(_02649_),
    .X(_02657_));
 sky130_fd_sc_hd__clkbuf_1 _19051_ (.A(_02657_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _19052_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.ready_buffer[57] ),
    .S(_02649_),
    .X(_02658_));
 sky130_fd_sc_hd__clkbuf_1 _19053_ (.A(_02658_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _19054_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.ready_buffer[58] ),
    .S(_02649_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_1 _19055_ (.A(_02659_),
    .X(_00691_));
 sky130_fd_sc_hd__buf_4 _19056_ (.A(_02593_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _19057_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _19058_ (.A(_02661_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _19059_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.ready_buffer[60] ),
    .S(_02660_),
    .X(_02662_));
 sky130_fd_sc_hd__clkbuf_1 _19060_ (.A(_02662_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _19061_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.ready_buffer[61] ),
    .S(_02660_),
    .X(_02663_));
 sky130_fd_sc_hd__clkbuf_1 _19062_ (.A(_02663_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _19063_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.ready_buffer[62] ),
    .S(_02660_),
    .X(_02664_));
 sky130_fd_sc_hd__clkbuf_1 _19064_ (.A(_02664_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _19065_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.ready_buffer[63] ),
    .S(_02660_),
    .X(_02665_));
 sky130_fd_sc_hd__clkbuf_1 _19066_ (.A(_02665_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _19067_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.ready_buffer[64] ),
    .S(_02660_),
    .X(_02666_));
 sky130_fd_sc_hd__clkbuf_1 _19068_ (.A(_02666_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _19069_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.ready_buffer[65] ),
    .S(_02660_),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _19070_ (.A(_02667_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _19071_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.ready_buffer[66] ),
    .S(_02660_),
    .X(_02668_));
 sky130_fd_sc_hd__clkbuf_1 _19072_ (.A(_02668_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _19073_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.ready_buffer[67] ),
    .S(_02660_),
    .X(_02669_));
 sky130_fd_sc_hd__clkbuf_1 _19074_ (.A(_02669_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _19075_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.ready_buffer[68] ),
    .S(_02660_),
    .X(_02670_));
 sky130_fd_sc_hd__clkbuf_1 _19076_ (.A(_02670_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _19077_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.ready_buffer[69] ),
    .S(_02594_),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_1 _19078_ (.A(_02671_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _19079_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.ready_buffer[70] ),
    .S(_02594_),
    .X(_02672_));
 sky130_fd_sc_hd__clkbuf_1 _19080_ (.A(_02672_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _19081_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.ready_buffer[71] ),
    .S(_02594_),
    .X(_02673_));
 sky130_fd_sc_hd__clkbuf_1 _19082_ (.A(_02673_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _19083_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.ready_buffer[72] ),
    .S(_02594_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_1 _19084_ (.A(_02674_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _19085_ (.A0(\rbzero.pov.spi_buffer[73] ),
    .A1(\rbzero.pov.ready_buffer[73] ),
    .S(_02594_),
    .X(_02675_));
 sky130_fd_sc_hd__clkbuf_1 _19086_ (.A(_02675_),
    .X(_00706_));
 sky130_fd_sc_hd__o311a_1 _19087_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(\rbzero.spi_registers.spi_counter[2] ),
    .A3(_02567_),
    .B1(_02558_),
    .C1(_02557_),
    .X(_02676_));
 sky130_fd_sc_hd__buf_4 _19088_ (.A(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _19089_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__clkbuf_1 _19090_ (.A(_02678_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _19091_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02677_),
    .X(_02679_));
 sky130_fd_sc_hd__clkbuf_1 _19092_ (.A(_02679_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _19093_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02677_),
    .X(_02680_));
 sky130_fd_sc_hd__clkbuf_1 _19094_ (.A(_02680_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _19095_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02677_),
    .X(_02681_));
 sky130_fd_sc_hd__clkbuf_1 _19096_ (.A(_02681_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _19097_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02677_),
    .X(_02682_));
 sky130_fd_sc_hd__clkbuf_1 _19098_ (.A(_02682_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _19099_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02677_),
    .X(_02683_));
 sky130_fd_sc_hd__clkbuf_1 _19100_ (.A(_02683_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _19101_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02677_),
    .X(_02684_));
 sky130_fd_sc_hd__clkbuf_1 _19102_ (.A(_02684_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _19103_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02677_),
    .X(_02685_));
 sky130_fd_sc_hd__clkbuf_1 _19104_ (.A(_02685_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _19105_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02677_),
    .X(_02686_));
 sky130_fd_sc_hd__clkbuf_1 _19106_ (.A(_02686_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _19107_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02677_),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_1 _19108_ (.A(_02687_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _19109_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02676_),
    .X(_02688_));
 sky130_fd_sc_hd__clkbuf_1 _19110_ (.A(_02688_),
    .X(_00717_));
 sky130_fd_sc_hd__nand2_1 _19111_ (.A(_02557_),
    .B(_02558_),
    .Y(_02689_));
 sky130_fd_sc_hd__or4_2 _19112_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .C(_02567_),
    .D(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _19113_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.spi_cmd[0] ),
    .S(_02690_),
    .X(_02691_));
 sky130_fd_sc_hd__clkbuf_1 _19114_ (.A(_02691_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _19115_ (.A0(\rbzero.spi_registers.spi_cmd[0] ),
    .A1(\rbzero.spi_registers.spi_cmd[1] ),
    .S(_02690_),
    .X(_02692_));
 sky130_fd_sc_hd__clkbuf_1 _19116_ (.A(_02692_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _19117_ (.A0(\rbzero.spi_registers.spi_cmd[1] ),
    .A1(\rbzero.spi_registers.spi_cmd[2] ),
    .S(_02690_),
    .X(_02693_));
 sky130_fd_sc_hd__clkbuf_1 _19118_ (.A(_02693_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _19119_ (.A0(\rbzero.spi_registers.spi_cmd[2] ),
    .A1(\rbzero.spi_registers.spi_cmd[3] ),
    .S(_02690_),
    .X(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _19120_ (.A(_02694_),
    .X(_00721_));
 sky130_fd_sc_hd__buf_6 _19121_ (.A(_03555_),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _19122_ (.A0(net42),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__clkbuf_1 _19123_ (.A(_02696_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _19124_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_05189_),
    .X(_02697_));
 sky130_fd_sc_hd__clkbuf_1 _19125_ (.A(_02697_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _19126_ (.A0(net41),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_02695_),
    .X(_02698_));
 sky130_fd_sc_hd__clkbuf_1 _19127_ (.A(_02698_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _19128_ (.A0(\rbzero.spi_registers.ss_buffer[1] ),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_05189_),
    .X(_02699_));
 sky130_fd_sc_hd__clkbuf_1 _19129_ (.A(_02699_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _19130_ (.A0(net43),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_02695_),
    .X(_02700_));
 sky130_fd_sc_hd__clkbuf_1 _19131_ (.A(_02700_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _19132_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_05189_),
    .X(_02701_));
 sky130_fd_sc_hd__clkbuf_1 _19133_ (.A(_02701_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _19134_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[2] ),
    .S(_02695_),
    .X(_02702_));
 sky130_fd_sc_hd__clkbuf_1 _19135_ (.A(_02702_),
    .X(_00728_));
 sky130_fd_sc_hd__nand3_2 _19136_ (.A(_04891_),
    .B(_04887_),
    .C(\gpout0.vpos[6] ),
    .Y(_02703_));
 sky130_fd_sc_hd__and3_1 _19137_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .X(_02704_));
 sky130_fd_sc_hd__and2_1 _19138_ (.A(\gpout0.vpos[3] ),
    .B(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__nand2_1 _19139_ (.A(_04037_),
    .B(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__nor4_4 _19140_ (.A(_04890_),
    .B(_04315_),
    .C(_02703_),
    .D(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__buf_4 _19141_ (.A(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__and2_1 _19142_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__buf_2 _19143_ (.A(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__clkbuf_4 _19144_ (.A(_02708_),
    .X(_02711_));
 sky130_fd_sc_hd__nand2_2 _19145_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__or2_1 _19146_ (.A(\rbzero.spi_registers.new_other[6] ),
    .B(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__clkbuf_4 _19147_ (.A(_05190_),
    .X(_02714_));
 sky130_fd_sc_hd__o211a_1 _19148_ (.A1(\rbzero.otherx[0] ),
    .A2(_02710_),
    .B1(_02713_),
    .C1(_02714_),
    .X(_00729_));
 sky130_fd_sc_hd__or2_1 _19149_ (.A(\rbzero.spi_registers.new_other[7] ),
    .B(_02712_),
    .X(_02715_));
 sky130_fd_sc_hd__o211a_1 _19150_ (.A1(\rbzero.otherx[1] ),
    .A2(_02710_),
    .B1(_02715_),
    .C1(_02714_),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _19151_ (.A(\rbzero.spi_registers.new_other[8] ),
    .B(_02712_),
    .X(_02716_));
 sky130_fd_sc_hd__o211a_1 _19152_ (.A1(\rbzero.otherx[2] ),
    .A2(_02710_),
    .B1(_02716_),
    .C1(_02714_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _19153_ (.A(\rbzero.spi_registers.new_other[9] ),
    .B(_02712_),
    .X(_02717_));
 sky130_fd_sc_hd__o211a_1 _19154_ (.A1(\rbzero.otherx[3] ),
    .A2(_02710_),
    .B1(_02717_),
    .C1(_02714_),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _19155_ (.A(\rbzero.spi_registers.new_other[10] ),
    .B(_02712_),
    .X(_02718_));
 sky130_fd_sc_hd__o211a_1 _19156_ (.A1(\rbzero.otherx[4] ),
    .A2(_02710_),
    .B1(_02718_),
    .C1(_02714_),
    .X(_00733_));
 sky130_fd_sc_hd__or2_1 _19157_ (.A(\rbzero.spi_registers.new_other[0] ),
    .B(_02712_),
    .X(_02719_));
 sky130_fd_sc_hd__o211a_1 _19158_ (.A1(\rbzero.othery[0] ),
    .A2(_02710_),
    .B1(_02719_),
    .C1(_02714_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _19159_ (.A(\rbzero.spi_registers.new_other[1] ),
    .B(_02712_),
    .X(_02720_));
 sky130_fd_sc_hd__buf_6 _19160_ (.A(_05189_),
    .X(_02721_));
 sky130_fd_sc_hd__buf_2 _19161_ (.A(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__o211a_1 _19162_ (.A1(\rbzero.othery[1] ),
    .A2(_02710_),
    .B1(_02720_),
    .C1(_02722_),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _19163_ (.A(\rbzero.spi_registers.new_other[2] ),
    .B(_02712_),
    .X(_02723_));
 sky130_fd_sc_hd__o211a_1 _19164_ (.A1(\rbzero.othery[2] ),
    .A2(_02710_),
    .B1(_02723_),
    .C1(_02722_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _19165_ (.A(\rbzero.spi_registers.new_other[3] ),
    .B(_02712_),
    .X(_02724_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(\rbzero.othery[3] ),
    .A2(_02710_),
    .B1(_02724_),
    .C1(_02722_),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _19167_ (.A(\rbzero.spi_registers.new_other[4] ),
    .B(_02712_),
    .X(_02725_));
 sky130_fd_sc_hd__o211a_1 _19168_ (.A1(\rbzero.othery[4] ),
    .A2(_02710_),
    .B1(_02725_),
    .C1(_02722_),
    .X(_00738_));
 sky130_fd_sc_hd__inv_2 _19169_ (.A(\rbzero.spi_registers.got_new_vinf ),
    .Y(_02726_));
 sky130_fd_sc_hd__or4_4 _19170_ (.A(\gpout0.vpos[9] ),
    .B(_04315_),
    .C(_02703_),
    .D(_02706_),
    .X(_02727_));
 sky130_fd_sc_hd__buf_4 _19171_ (.A(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__a21o_1 _19172_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_02711_),
    .B1(\rbzero.row_render.vinf ),
    .X(_02729_));
 sky130_fd_sc_hd__buf_4 _19173_ (.A(_05190_),
    .X(_02730_));
 sky130_fd_sc_hd__o311a_1 _19174_ (.A1(\rbzero.spi_registers.new_vinf ),
    .A2(_02726_),
    .A3(_02728_),
    .B1(_02729_),
    .C1(_02730_),
    .X(_00739_));
 sky130_fd_sc_hd__and2_1 _19175_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02708_),
    .X(_02731_));
 sky130_fd_sc_hd__clkbuf_2 _19176_ (.A(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__nand2_1 _19177_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02711_),
    .Y(_02733_));
 sky130_fd_sc_hd__or2_1 _19178_ (.A(\rbzero.spi_registers.new_leak[0] ),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__o211a_1 _19179_ (.A1(\rbzero.floor_leak[0] ),
    .A2(_02732_),
    .B1(_02734_),
    .C1(_02722_),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _19180_ (.A(\rbzero.spi_registers.new_leak[1] ),
    .B(_02733_),
    .X(_02735_));
 sky130_fd_sc_hd__o211a_1 _19181_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_02732_),
    .B1(_02735_),
    .C1(_02722_),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _19182_ (.A(\rbzero.spi_registers.new_leak[2] ),
    .B(_02733_),
    .X(_02736_));
 sky130_fd_sc_hd__o211a_1 _19183_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_02732_),
    .B1(_02736_),
    .C1(_02722_),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _19184_ (.A(\rbzero.spi_registers.new_leak[3] ),
    .B(_02733_),
    .X(_02737_));
 sky130_fd_sc_hd__o211a_1 _19185_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_02732_),
    .B1(_02737_),
    .C1(_02722_),
    .X(_00743_));
 sky130_fd_sc_hd__or2_1 _19186_ (.A(\rbzero.spi_registers.new_leak[4] ),
    .B(_02733_),
    .X(_02738_));
 sky130_fd_sc_hd__o211a_1 _19187_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_02732_),
    .B1(_02738_),
    .C1(_02722_),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _19188_ (.A(\rbzero.spi_registers.new_leak[5] ),
    .B(_02733_),
    .X(_02739_));
 sky130_fd_sc_hd__o211a_1 _19189_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_02732_),
    .B1(_02739_),
    .C1(_02722_),
    .X(_00745_));
 sky130_fd_sc_hd__nand2_2 _19190_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_02707_),
    .Y(_02740_));
 sky130_fd_sc_hd__buf_6 _19191_ (.A(_03555_),
    .X(_02741_));
 sky130_fd_sc_hd__a31o_1 _19192_ (.A1(\rbzero.spi_registers.new_sky[0] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02711_),
    .B1(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__a21o_1 _19193_ (.A1(\rbzero.color_sky[0] ),
    .A2(_02740_),
    .B1(_02742_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _19194_ (.A0(\rbzero.spi_registers.new_sky[1] ),
    .A1(\rbzero.color_sky[1] ),
    .S(_02740_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_1 _19195_ (.A(_09753_),
    .B(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_1 _19196_ (.A(_02744_),
    .X(_00747_));
 sky130_fd_sc_hd__a31o_1 _19197_ (.A1(\rbzero.spi_registers.new_sky[2] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02711_),
    .B1(_02741_),
    .X(_02745_));
 sky130_fd_sc_hd__a21o_1 _19198_ (.A1(\rbzero.color_sky[2] ),
    .A2(_02740_),
    .B1(_02745_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _19199_ (.A0(\rbzero.spi_registers.new_sky[3] ),
    .A1(\rbzero.color_sky[3] ),
    .S(_02740_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_1 _19200_ (.A(_09753_),
    .B(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__clkbuf_1 _19201_ (.A(_02747_),
    .X(_00749_));
 sky130_fd_sc_hd__a31o_1 _19202_ (.A1(\rbzero.spi_registers.new_sky[4] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02711_),
    .B1(_02741_),
    .X(_02748_));
 sky130_fd_sc_hd__a21o_1 _19203_ (.A1(\rbzero.color_sky[4] ),
    .A2(_02740_),
    .B1(_02748_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _19204_ (.A0(\rbzero.spi_registers.new_sky[5] ),
    .A1(\rbzero.color_sky[5] ),
    .S(_02740_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_1 _19205_ (.A(_09753_),
    .B(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__clkbuf_1 _19206_ (.A(_02750_),
    .X(_00751_));
 sky130_fd_sc_hd__nand2_2 _19207_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_02707_),
    .Y(_02751_));
 sky130_fd_sc_hd__mux2_1 _19208_ (.A0(\rbzero.spi_registers.new_floor[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_1 _19209_ (.A(_09753_),
    .B(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__clkbuf_1 _19210_ (.A(_02753_),
    .X(_00752_));
 sky130_fd_sc_hd__a31o_1 _19211_ (.A1(\rbzero.spi_registers.new_floor[1] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02711_),
    .B1(_03911_),
    .X(_02754_));
 sky130_fd_sc_hd__a21o_1 _19212_ (.A1(\rbzero.color_floor[1] ),
    .A2(_02751_),
    .B1(_02754_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _19213_ (.A0(\rbzero.spi_registers.new_floor[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_02751_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_1 _19214_ (.A(_09753_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__clkbuf_1 _19215_ (.A(_02756_),
    .X(_00754_));
 sky130_fd_sc_hd__a31o_1 _19216_ (.A1(\rbzero.spi_registers.new_floor[3] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02711_),
    .B1(_03911_),
    .X(_02757_));
 sky130_fd_sc_hd__a21o_1 _19217_ (.A1(\rbzero.color_floor[3] ),
    .A2(_02751_),
    .B1(_02757_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _19218_ (.A0(\rbzero.spi_registers.new_floor[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_02751_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_1 _19219_ (.A(_09753_),
    .B(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__clkbuf_1 _19220_ (.A(_02759_),
    .X(_00756_));
 sky130_fd_sc_hd__a31o_1 _19221_ (.A1(\rbzero.spi_registers.new_floor[5] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02711_),
    .B1(_03911_),
    .X(_02760_));
 sky130_fd_sc_hd__a21o_1 _19222_ (.A1(\rbzero.color_floor[5] ),
    .A2(_02751_),
    .B1(_02760_),
    .X(_00757_));
 sky130_fd_sc_hd__and2_1 _19223_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02708_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_2 _19224_ (.A(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__nand2_2 _19225_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02711_),
    .Y(_02763_));
 sky130_fd_sc_hd__or2_1 _19226_ (.A(\rbzero.spi_registers.new_vshift[0] ),
    .B(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__buf_4 _19227_ (.A(_02721_),
    .X(_02765_));
 sky130_fd_sc_hd__o211a_1 _19228_ (.A1(\rbzero.spi_registers.vshift[0] ),
    .A2(_02762_),
    .B1(_02764_),
    .C1(_02765_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _19229_ (.A(\rbzero.spi_registers.new_vshift[1] ),
    .B(_02763_),
    .X(_02766_));
 sky130_fd_sc_hd__o211a_1 _19230_ (.A1(\rbzero.spi_registers.vshift[1] ),
    .A2(_02762_),
    .B1(_02766_),
    .C1(_02765_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _19231_ (.A(\rbzero.spi_registers.new_vshift[2] ),
    .B(_02763_),
    .X(_02767_));
 sky130_fd_sc_hd__o211a_1 _19232_ (.A1(\rbzero.spi_registers.vshift[2] ),
    .A2(_02762_),
    .B1(_02767_),
    .C1(_02765_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _19233_ (.A(\rbzero.spi_registers.new_vshift[3] ),
    .B(_02763_),
    .X(_02768_));
 sky130_fd_sc_hd__o211a_1 _19234_ (.A1(\rbzero.spi_registers.vshift[3] ),
    .A2(_02762_),
    .B1(_02768_),
    .C1(_02765_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19235_ (.A(\rbzero.spi_registers.new_vshift[4] ),
    .B(_02763_),
    .X(_02769_));
 sky130_fd_sc_hd__o211a_1 _19236_ (.A1(\rbzero.spi_registers.vshift[4] ),
    .A2(_02762_),
    .B1(_02769_),
    .C1(_02765_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19237_ (.A(\rbzero.spi_registers.new_vshift[5] ),
    .B(_02763_),
    .X(_02770_));
 sky130_fd_sc_hd__o211a_1 _19238_ (.A1(\rbzero.spi_registers.vshift[5] ),
    .A2(_02762_),
    .B1(_02770_),
    .C1(_02765_),
    .X(_00763_));
 sky130_fd_sc_hd__and4b_1 _19239_ (.A_N(\rbzero.spi_registers.spi_done ),
    .B(_02557_),
    .C(_02558_),
    .D(_02572_),
    .X(_02771_));
 sky130_fd_sc_hd__clkbuf_1 _19240_ (.A(_02771_),
    .X(_00764_));
 sky130_fd_sc_hd__nand3_1 _19241_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_03480_),
    .C(_02560_),
    .Y(_02772_));
 sky130_fd_sc_hd__or2_1 _19242_ (.A(_02561_),
    .B(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__clkbuf_4 _19243_ (.A(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _19244_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__clkbuf_1 _19245_ (.A(_02775_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _19246_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_02774_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _19247_ (.A(_02776_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _19248_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_02774_),
    .X(_02777_));
 sky130_fd_sc_hd__clkbuf_1 _19249_ (.A(_02777_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _19250_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_02774_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _19251_ (.A(_02778_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _19252_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_02774_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_1 _19253_ (.A(_02779_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _19254_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_02774_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_1 _19255_ (.A(_02780_),
    .X(_00770_));
 sky130_fd_sc_hd__inv_2 _19256_ (.A(_02774_),
    .Y(_02781_));
 sky130_fd_sc_hd__a31o_1 _19257_ (.A1(\rbzero.spi_registers.got_new_sky ),
    .A2(_02730_),
    .A3(_02728_),
    .B1(_02781_),
    .X(_00771_));
 sky130_fd_sc_hd__or3b_1 _19258_ (.A(_02772_),
    .B(\rbzero.spi_registers.spi_cmd[1] ),
    .C_N(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_4 _19259_ (.A(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _19260_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_floor[0] ),
    .S(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _19261_ (.A(_02784_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _19262_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_floor[1] ),
    .S(_02783_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_1 _19263_ (.A(_02785_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _19264_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_floor[2] ),
    .S(_02783_),
    .X(_02786_));
 sky130_fd_sc_hd__clkbuf_1 _19265_ (.A(_02786_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _19266_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_floor[3] ),
    .S(_02783_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_1 _19267_ (.A(_02787_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _19268_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_floor[4] ),
    .S(_02783_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _19269_ (.A(_02788_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _19270_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_floor[5] ),
    .S(_02783_),
    .X(_02789_));
 sky130_fd_sc_hd__clkbuf_1 _19271_ (.A(_02789_),
    .X(_00777_));
 sky130_fd_sc_hd__inv_2 _19272_ (.A(_02783_),
    .Y(_02790_));
 sky130_fd_sc_hd__a31o_1 _19273_ (.A1(\rbzero.spi_registers.got_new_floor ),
    .A2(_02730_),
    .A3(_02728_),
    .B1(_02790_),
    .X(_00778_));
 sky130_fd_sc_hd__or3b_1 _19274_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02772_),
    .C_N(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_4 _19275_ (.A(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _19276_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.new_leak[0] ),
    .S(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__clkbuf_1 _19277_ (.A(_02793_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _19278_ (.A0(\rbzero.spi_registers.spi_buffer[1] ),
    .A1(\rbzero.spi_registers.new_leak[1] ),
    .S(_02792_),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_1 _19279_ (.A(_02794_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _19280_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.new_leak[2] ),
    .S(_02792_),
    .X(_02795_));
 sky130_fd_sc_hd__clkbuf_1 _19281_ (.A(_02795_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _19282_ (.A0(\rbzero.spi_registers.spi_buffer[3] ),
    .A1(\rbzero.spi_registers.new_leak[3] ),
    .S(_02792_),
    .X(_02796_));
 sky130_fd_sc_hd__clkbuf_1 _19283_ (.A(_02796_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _19284_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.new_leak[4] ),
    .S(_02792_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_1 _19285_ (.A(_02797_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _19286_ (.A0(\rbzero.spi_registers.spi_buffer[5] ),
    .A1(\rbzero.spi_registers.new_leak[5] ),
    .S(_02792_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _19287_ (.A(_02798_),
    .X(_00784_));
 sky130_fd_sc_hd__inv_2 _19288_ (.A(_02792_),
    .Y(_02799_));
 sky130_fd_sc_hd__a31o_1 _19289_ (.A1(\rbzero.spi_registers.got_new_leak ),
    .A2(_02730_),
    .A3(_02728_),
    .B1(_02799_),
    .X(_00785_));
 sky130_fd_sc_hd__and3_1 _19290_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_03480_),
    .C(_02569_),
    .X(_02800_));
 sky130_fd_sc_hd__buf_4 _19291_ (.A(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _19292_ (.A0(\rbzero.spi_registers.new_other[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_1 _19293_ (.A(_02802_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _19294_ (.A0(\rbzero.spi_registers.new_other[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02801_),
    .X(_02803_));
 sky130_fd_sc_hd__clkbuf_1 _19295_ (.A(_02803_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _19296_ (.A0(\rbzero.spi_registers.new_other[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02801_),
    .X(_02804_));
 sky130_fd_sc_hd__clkbuf_1 _19297_ (.A(_02804_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _19298_ (.A0(\rbzero.spi_registers.new_other[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02801_),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_1 _19299_ (.A(_02805_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _19300_ (.A0(\rbzero.spi_registers.new_other[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02801_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _19301_ (.A(_02806_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _19302_ (.A0(\rbzero.spi_registers.new_other[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02801_),
    .X(_02807_));
 sky130_fd_sc_hd__clkbuf_1 _19303_ (.A(_02807_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _19304_ (.A0(\rbzero.spi_registers.new_other[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02801_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _19305_ (.A(_02808_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _19306_ (.A0(\rbzero.spi_registers.new_other[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02801_),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _19307_ (.A(_02809_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _19308_ (.A0(\rbzero.spi_registers.new_other[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02801_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_1 _19309_ (.A(_02810_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _19310_ (.A0(\rbzero.spi_registers.new_other[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02800_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_1 _19311_ (.A(_02811_),
    .X(_00795_));
 sky130_fd_sc_hd__a31o_1 _19312_ (.A1(\rbzero.spi_registers.got_new_other ),
    .A2(_02730_),
    .A3(_02728_),
    .B1(_02801_),
    .X(_00796_));
 sky130_fd_sc_hd__and3_1 _19313_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_03480_),
    .C(_02563_),
    .X(_02812_));
 sky130_fd_sc_hd__clkbuf_4 _19314_ (.A(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _19315_ (.A0(\rbzero.spi_registers.new_vshift[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__clkbuf_1 _19316_ (.A(_02814_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _19317_ (.A0(\rbzero.spi_registers.new_vshift[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02813_),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_1 _19318_ (.A(_02815_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _19319_ (.A0(\rbzero.spi_registers.new_vshift[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_02813_),
    .X(_02816_));
 sky130_fd_sc_hd__clkbuf_1 _19320_ (.A(_02816_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _19321_ (.A0(\rbzero.spi_registers.new_vshift[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02813_),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _19322_ (.A(_02817_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _19323_ (.A0(\rbzero.spi_registers.new_vshift[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_02813_),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_1 _19324_ (.A(_02818_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _19325_ (.A0(\rbzero.spi_registers.new_vshift[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02813_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _19326_ (.A(_02819_),
    .X(_00802_));
 sky130_fd_sc_hd__a31o_1 _19327_ (.A1(\rbzero.spi_registers.got_new_vshift ),
    .A2(_02730_),
    .A3(_02728_),
    .B1(_02813_),
    .X(_00803_));
 sky130_fd_sc_hd__nor2_4 _19328_ (.A(net39),
    .B(net38),
    .Y(_02820_));
 sky130_fd_sc_hd__or2_1 _19329_ (.A(_02728_),
    .B(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_4 _19330_ (.A(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__clkbuf_4 _19331_ (.A(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__o211a_1 _19332_ (.A1(\rbzero.pov.spi_done ),
    .A2(\rbzero.pov.ready ),
    .B1(_02730_),
    .C1(_02823_),
    .X(_00804_));
 sky130_fd_sc_hd__nor2_1 _19333_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_1 _19334_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02825_));
 sky130_fd_sc_hd__and2b_1 _19335_ (.A_N(_02824_),
    .B(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__or2_1 _19336_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .X(_02827_));
 sky130_fd_sc_hd__nor2_1 _19337_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02828_));
 sky130_fd_sc_hd__nand2_1 _19338_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _19339_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .Y(_02830_));
 sky130_fd_sc_hd__or2_1 _19340_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_02831_));
 sky130_fd_sc_hd__nand3b_1 _19341_ (.A_N(_02830_),
    .B(_02831_),
    .C(_02829_),
    .Y(_02832_));
 sky130_fd_sc_hd__and2_1 _19342_ (.A(_02829_),
    .B(_02832_),
    .X(_02833_));
 sky130_fd_sc_hd__nand2_1 _19343_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02834_));
 sky130_fd_sc_hd__o21ai_1 _19344_ (.A1(_02828_),
    .A2(_02833_),
    .B1(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _19345_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_02836_));
 sky130_fd_sc_hd__a21boi_1 _19346_ (.A1(_02827_),
    .A2(_02835_),
    .B1_N(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__xnor2_1 _19347_ (.A(_02826_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a22o_1 _19348_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_07703_),
    .B1(_07855_),
    .B2(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_02839_));
 sky130_fd_sc_hd__a21o_1 _19349_ (.A1(_07728_),
    .A2(_02838_),
    .B1(_02839_),
    .X(_00805_));
 sky130_fd_sc_hd__nor2_1 _19350_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_02840_));
 sky130_fd_sc_hd__and2_1 _19351_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02841_));
 sky130_fd_sc_hd__o21ai_1 _19352_ (.A1(_02824_),
    .A2(_02837_),
    .B1(_02825_),
    .Y(_02842_));
 sky130_fd_sc_hd__or3_1 _19353_ (.A(_02840_),
    .B(_02841_),
    .C(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__o21ai_1 _19354_ (.A1(_02840_),
    .A2(_02841_),
    .B1(_02842_),
    .Y(_02844_));
 sky130_fd_sc_hd__a21oi_1 _19355_ (.A1(_02843_),
    .A2(_02844_),
    .B1(_07703_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _19356_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02846_));
 sky130_fd_sc_hd__or2_1 _19357_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_02847_));
 sky130_fd_sc_hd__a31o_1 _19358_ (.A1(_07703_),
    .A2(_02846_),
    .A3(_02847_),
    .B1(_07706_),
    .X(_02848_));
 sky130_fd_sc_hd__o22a_1 _19359_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_00013_),
    .B1(_02845_),
    .B2(_02848_),
    .X(_00806_));
 sky130_fd_sc_hd__or2_1 _19360_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02847_),
    .X(_02849_));
 sky130_fd_sc_hd__nand2_1 _19361_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02847_),
    .Y(_02850_));
 sky130_fd_sc_hd__nor2_1 _19362_ (.A(_04471_),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02851_));
 sky130_fd_sc_hd__nand2_1 _19363_ (.A(_04471_),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02852_));
 sky130_fd_sc_hd__or2b_1 _19364_ (.A(_02851_),
    .B_N(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__or2_1 _19365_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02854_));
 sky130_fd_sc_hd__a21oi_1 _19366_ (.A1(_02854_),
    .A2(_02842_),
    .B1(_02841_),
    .Y(_02855_));
 sky130_fd_sc_hd__xnor2_1 _19367_ (.A(_02853_),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__nor2_1 _19368_ (.A(_07676_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__a31o_1 _19369_ (.A1(_07676_),
    .A2(_02849_),
    .A3(_02850_),
    .B1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__mux2_1 _19370_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(_02858_),
    .S(_07718_),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _19371_ (.A(_02859_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _19372_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02860_));
 sky130_fd_sc_hd__nand2_1 _19373_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_02861_));
 sky130_fd_sc_hd__nand2_1 _19374_ (.A(_02860_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__o21ai_1 _19375_ (.A1(_02851_),
    .A2(_02855_),
    .B1(_02852_),
    .Y(_02863_));
 sky130_fd_sc_hd__xnor2_1 _19376_ (.A(_02862_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__or2_1 _19377_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_02849_),
    .X(_02865_));
 sky130_fd_sc_hd__a21oi_1 _19378_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(_02849_),
    .B1(_04034_),
    .Y(_02866_));
 sky130_fd_sc_hd__a221o_1 _19379_ (.A1(_04034_),
    .A2(_02864_),
    .B1(_02865_),
    .B2(_02866_),
    .C1(_07706_),
    .X(_02867_));
 sky130_fd_sc_hd__o21a_1 _19380_ (.A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A2(_00013_),
    .B1(_02867_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19381_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02868_));
 sky130_fd_sc_hd__nand2_1 _19382_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_02869_));
 sky130_fd_sc_hd__nand2_1 _19383_ (.A(_02868_),
    .B(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__a21bo_1 _19384_ (.A1(_02860_),
    .A2(_02863_),
    .B1_N(_02861_),
    .X(_02871_));
 sky130_fd_sc_hd__xnor2_1 _19385_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__or2_1 _19386_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_02873_));
 sky130_fd_sc_hd__nand2_1 _19387_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02874_));
 sky130_fd_sc_hd__nand2_1 _19388_ (.A(_02873_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__xnor2_1 _19389_ (.A(_02865_),
    .B(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__a22o_1 _19390_ (.A1(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2(_07706_),
    .B1(_02876_),
    .B2(_07703_),
    .X(_02877_));
 sky130_fd_sc_hd__a21o_1 _19391_ (.A1(_07728_),
    .A2(_02872_),
    .B1(_02877_),
    .X(_00809_));
 sky130_fd_sc_hd__a21bo_1 _19392_ (.A1(_02868_),
    .A2(_02871_),
    .B1_N(_02869_),
    .X(_02878_));
 sky130_fd_sc_hd__or2_1 _19393_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02879_));
 sky130_fd_sc_hd__nand2_1 _19394_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_02880_));
 sky130_fd_sc_hd__nand2_1 _19395_ (.A(_02879_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__xnor2_1 _19396_ (.A(_02878_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_1 _19397_ (.A(_02865_),
    .B(_02875_),
    .Y(_02883_));
 sky130_fd_sc_hd__and2_1 _19398_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_02884_));
 sky130_fd_sc_hd__nor2_1 _19399_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_02885_));
 sky130_fd_sc_hd__o21ai_1 _19400_ (.A1(_02884_),
    .A2(_02885_),
    .B1(_02873_),
    .Y(_02886_));
 sky130_fd_sc_hd__or3_1 _19401_ (.A(_02873_),
    .B(_02884_),
    .C(_02885_),
    .X(_02887_));
 sky130_fd_sc_hd__and2_1 _19402_ (.A(_02886_),
    .B(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__or2_1 _19403_ (.A(_02883_),
    .B(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_1 _19404_ (.A(_02883_),
    .B(_02888_),
    .Y(_02890_));
 sky130_fd_sc_hd__a31o_1 _19405_ (.A1(_03913_),
    .A2(_02889_),
    .A3(_02890_),
    .B1(_07695_),
    .X(_02891_));
 sky130_fd_sc_hd__a21o_1 _19406_ (.A1(_04035_),
    .A2(_02882_),
    .B1(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__o21a_1 _19407_ (.A1(\rbzero.wall_tracer.rayAddendY[0] ),
    .A2(_00013_),
    .B1(_02892_),
    .X(_00810_));
 sky130_fd_sc_hd__nand2_1 _19408_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_02893_));
 sky130_fd_sc_hd__or2_1 _19409_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02894_));
 sky130_fd_sc_hd__or2b_1 _19410_ (.A(_02878_),
    .B_N(_02880_),
    .X(_02895_));
 sky130_fd_sc_hd__nand4_2 _19411_ (.A(_02879_),
    .B(_02893_),
    .C(_02894_),
    .D(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__a22o_1 _19412_ (.A1(_02893_),
    .A2(_02894_),
    .B1(_02895_),
    .B2(_02879_),
    .X(_02897_));
 sky130_fd_sc_hd__xnor2_1 _19413_ (.A(_04471_),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_02898_));
 sky130_fd_sc_hd__a21o_1 _19414_ (.A1(_02887_),
    .A2(_02890_),
    .B1(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__nand3_1 _19415_ (.A(_02887_),
    .B(_02890_),
    .C(_02898_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _19416_ (.A(_02899_),
    .B(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__xnor2_1 _19417_ (.A(_02885_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__a22o_1 _19418_ (.A1(\rbzero.wall_tracer.rayAddendY[1] ),
    .A2(_07695_),
    .B1(_02902_),
    .B2(_07703_),
    .X(_02903_));
 sky130_fd_sc_hd__a31o_1 _19419_ (.A1(_07756_),
    .A2(_02896_),
    .A3(_02897_),
    .B1(_02903_),
    .X(_00811_));
 sky130_fd_sc_hd__clkbuf_4 _19420_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_02904_));
 sky130_fd_sc_hd__buf_2 _19421_ (.A(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__buf_4 _19422_ (.A(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__xnor2_1 _19423_ (.A(_02906_),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_02907_));
 sky130_fd_sc_hd__a21oi_1 _19424_ (.A1(_02893_),
    .A2(_02896_),
    .B1(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__a31o_1 _19425_ (.A1(_02893_),
    .A2(_02896_),
    .A3(_02907_),
    .B1(_07676_),
    .X(_02909_));
 sky130_fd_sc_hd__and2_1 _19426_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_02910_));
 sky130_fd_sc_hd__nor2_1 _19427_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .Y(_02911_));
 sky130_fd_sc_hd__o22ai_1 _19428_ (.A1(_04471_),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .B1(_02910_),
    .B2(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__or4_1 _19429_ (.A(_04471_),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .C(_02910_),
    .D(_02911_),
    .X(_02913_));
 sky130_fd_sc_hd__nand2_1 _19430_ (.A(_02912_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__a21bo_1 _19431_ (.A1(_02890_),
    .A2(_02898_),
    .B1_N(_02885_),
    .X(_02915_));
 sky130_fd_sc_hd__a21o_1 _19432_ (.A1(_02899_),
    .A2(_02915_),
    .B1(_02914_),
    .X(_02916_));
 sky130_fd_sc_hd__nand2_1 _19433_ (.A(_03912_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a31o_1 _19434_ (.A1(_02899_),
    .A2(_02914_),
    .A3(_02915_),
    .B1(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__o21ai_1 _19435_ (.A1(_02908_),
    .A2(_02909_),
    .B1(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__mux2_1 _19436_ (.A0(\rbzero.wall_tracer.rayAddendY[2] ),
    .A1(_02919_),
    .S(_07718_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _19437_ (.A(_02920_),
    .X(_00812_));
 sky130_fd_sc_hd__o21ai_1 _19438_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(\rbzero.debug_overlay.vplaneY[10] ),
    .Y(_02921_));
 sky130_fd_sc_hd__o21bai_1 _19439_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1_N(_02896_),
    .Y(_02922_));
 sky130_fd_sc_hd__and2_1 _19440_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02923_));
 sky130_fd_sc_hd__nor2_1 _19441_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02924_));
 sky130_fd_sc_hd__a211oi_2 _19442_ (.A1(_02921_),
    .A2(_02922_),
    .B1(_02923_),
    .C1(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__o211a_1 _19443_ (.A1(_02923_),
    .A2(_02924_),
    .B1(_02921_),
    .C1(_02922_),
    .X(_02926_));
 sky130_fd_sc_hd__or2_1 _19444_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_02927_));
 sky130_fd_sc_hd__nand2_1 _19445_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_1 _19446_ (.A(_02927_),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__a21oi_1 _19447_ (.A1(_02913_),
    .A2(_02916_),
    .B1(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__and3_1 _19448_ (.A(_02913_),
    .B(_02916_),
    .C(_02929_),
    .X(_02931_));
 sky130_fd_sc_hd__o21bai_1 _19449_ (.A1(_02930_),
    .A2(_02931_),
    .B1_N(_02911_),
    .Y(_02932_));
 sky130_fd_sc_hd__o41a_1 _19450_ (.A1(\rbzero.debug_overlay.vplaneY[-2] ),
    .A2(\rbzero.debug_overlay.vplaneY[-6] ),
    .A3(_02930_),
    .A4(_02931_),
    .B1(_03913_),
    .X(_02933_));
 sky130_fd_sc_hd__a22oi_1 _19451_ (.A1(\rbzero.wall_tracer.rayAddendY[3] ),
    .A2(_07855_),
    .B1(_02932_),
    .B2(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__o31ai_1 _19452_ (.A1(_07831_),
    .A2(_02925_),
    .A3(_02926_),
    .B1(_02934_),
    .Y(_00813_));
 sky130_fd_sc_hd__xor2_1 _19453_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_02935_));
 sky130_fd_sc_hd__or3_1 _19454_ (.A(_02923_),
    .B(_02925_),
    .C(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__o21ai_1 _19455_ (.A1(_02923_),
    .A2(_02925_),
    .B1(_02935_),
    .Y(_02937_));
 sky130_fd_sc_hd__nor2_1 _19456_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .Y(_02938_));
 sky130_fd_sc_hd__and2_1 _19457_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_02939_));
 sky130_fd_sc_hd__o21a_1 _19458_ (.A1(_02938_),
    .A2(_02939_),
    .B1(_02927_),
    .X(_02940_));
 sky130_fd_sc_hd__nor3_1 _19459_ (.A(_02927_),
    .B(_02938_),
    .C(_02939_),
    .Y(_02941_));
 sky130_fd_sc_hd__nor2_1 _19460_ (.A(_02940_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__o2bb2a_1 _19461_ (.A1_N(_02916_),
    .A2_N(_02929_),
    .B1(_02930_),
    .B2(_02911_),
    .X(_02943_));
 sky130_fd_sc_hd__and2_1 _19462_ (.A(_02942_),
    .B(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__o21ai_1 _19463_ (.A1(_02942_),
    .A2(_02943_),
    .B1(_07676_),
    .Y(_02945_));
 sky130_fd_sc_hd__o21ai_1 _19464_ (.A1(_02944_),
    .A2(_02945_),
    .B1(_04029_),
    .Y(_02946_));
 sky130_fd_sc_hd__a31o_1 _19465_ (.A1(_04035_),
    .A2(_02936_),
    .A3(_02937_),
    .B1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__o21a_1 _19466_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(_00013_),
    .B1(_02947_),
    .X(_00814_));
 sky130_fd_sc_hd__nand2_1 _19467_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_02948_));
 sky130_fd_sc_hd__or2_1 _19468_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_02949_));
 sky130_fd_sc_hd__nand2_1 _19469_ (.A(_02948_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__nand2_1 _19470_ (.A(_02925_),
    .B(_02935_),
    .Y(_02951_));
 sky130_fd_sc_hd__o21ai_2 _19471_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02904_),
    .Y(_02952_));
 sky130_fd_sc_hd__nand3_1 _19472_ (.A(_02950_),
    .B(_02951_),
    .C(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__a21o_1 _19473_ (.A1(_02951_),
    .A2(_02952_),
    .B1(_02950_),
    .X(_02954_));
 sky130_fd_sc_hd__and3_1 _19474_ (.A(_07678_),
    .B(_02953_),
    .C(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__xor2_1 _19475_ (.A(_02904_),
    .B(_04471_),
    .X(_02956_));
 sky130_fd_sc_hd__xor2_1 _19476_ (.A(_02938_),
    .B(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__o21a_1 _19477_ (.A1(_02941_),
    .A2(_02944_),
    .B1(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__nor2_1 _19478_ (.A(_04034_),
    .B(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__o31a_1 _19479_ (.A1(_02941_),
    .A2(_02944_),
    .A3(_02957_),
    .B1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__a211o_1 _19480_ (.A1(\rbzero.wall_tracer.rayAddendY[5] ),
    .A2(_07855_),
    .B1(_02955_),
    .C1(_02960_),
    .X(_00815_));
 sky130_fd_sc_hd__nor2_1 _19481_ (.A(_02905_),
    .B(\rbzero.debug_overlay.vplaneY[-2] ),
    .Y(_02961_));
 sky130_fd_sc_hd__and2_1 _19482_ (.A(_02905_),
    .B(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_02962_));
 sky130_fd_sc_hd__o22ai_1 _19483_ (.A1(_02905_),
    .A2(_04471_),
    .B1(_02961_),
    .B2(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__or3b_1 _19484_ (.A(_02905_),
    .B(_04471_),
    .C_N(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_02964_));
 sky130_fd_sc_hd__nand2_1 _19485_ (.A(_02963_),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__a21o_1 _19486_ (.A1(_02938_),
    .A2(_02956_),
    .B1(_02958_),
    .X(_02966_));
 sky130_fd_sc_hd__xnor2_1 _19487_ (.A(_02965_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__xor2_1 _19488_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_02968_));
 sky130_fd_sc_hd__nand2_1 _19489_ (.A(_02948_),
    .B(_02954_),
    .Y(_02969_));
 sky130_fd_sc_hd__xor2_1 _19490_ (.A(_02968_),
    .B(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _19491_ (.A0(_02967_),
    .A1(_02970_),
    .S(_04033_),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _19492_ (.A0(\rbzero.wall_tracer.rayAddendY[6] ),
    .A1(_02971_),
    .S(_07718_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _19493_ (.A(_02972_),
    .X(_00816_));
 sky130_fd_sc_hd__nand2_1 _19494_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_02973_));
 sky130_fd_sc_hd__or2_1 _19495_ (.A(_02904_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02974_));
 sky130_fd_sc_hd__nand2_1 _19496_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__or3b_1 _19497_ (.A(_02950_),
    .B(_02951_),
    .C_N(_02968_),
    .X(_02976_));
 sky130_fd_sc_hd__o21ai_1 _19498_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .B1(_02905_),
    .Y(_02977_));
 sky130_fd_sc_hd__nand4_1 _19499_ (.A(_02952_),
    .B(_02975_),
    .C(_02976_),
    .D(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__a31o_1 _19500_ (.A1(_02952_),
    .A2(_02976_),
    .A3(_02977_),
    .B1(_02975_),
    .X(_02979_));
 sky130_fd_sc_hd__or2_1 _19501_ (.A(_02905_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_02980_));
 sky130_fd_sc_hd__nand2_1 _19502_ (.A(_02905_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_02981_));
 sky130_fd_sc_hd__a21o_1 _19503_ (.A1(_02980_),
    .A2(_02981_),
    .B1(_02961_),
    .X(_02982_));
 sky130_fd_sc_hd__nand2_1 _19504_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_02961_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_1 _19505_ (.A(_02982_),
    .B(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__a21boi_1 _19506_ (.A1(_02963_),
    .A2(_02966_),
    .B1_N(_02964_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2_1 _19507_ (.A(_02984_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__or2_1 _19508_ (.A(_02984_),
    .B(_02985_),
    .X(_02987_));
 sky130_fd_sc_hd__a32o_1 _19509_ (.A1(_03913_),
    .A2(_02986_),
    .A3(_02987_),
    .B1(_07855_),
    .B2(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02988_));
 sky130_fd_sc_hd__a31o_1 _19510_ (.A1(_07679_),
    .A2(_02978_),
    .A3(_02979_),
    .B1(_02988_),
    .X(_00817_));
 sky130_fd_sc_hd__xnor2_1 _19511_ (.A(_02905_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_02989_));
 sky130_fd_sc_hd__a21oi_1 _19512_ (.A1(_02973_),
    .A2(_02979_),
    .B1(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__a31o_1 _19513_ (.A1(_02973_),
    .A2(_02979_),
    .A3(_02989_),
    .B1(_03913_),
    .X(_02991_));
 sky130_fd_sc_hd__nor2_1 _19514_ (.A(_02990_),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__and2_1 _19515_ (.A(_02906_),
    .B(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_02993_));
 sky130_fd_sc_hd__or2_1 _19516_ (.A(_02905_),
    .B(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_1 _19517_ (.A(_02980_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__o22a_1 _19518_ (.A1(\rbzero.debug_overlay.vplaneY[0] ),
    .A2(_02980_),
    .B1(_02993_),
    .B2(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__nand3_1 _19519_ (.A(_02983_),
    .B(_02987_),
    .C(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21o_1 _19520_ (.A1(_02983_),
    .A2(_02987_),
    .B1(_02996_),
    .X(_02998_));
 sky130_fd_sc_hd__a31o_1 _19521_ (.A1(_03913_),
    .A2(_02997_),
    .A3(_02998_),
    .B1(_07695_),
    .X(_02999_));
 sky130_fd_sc_hd__o22a_1 _19522_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(_00013_),
    .B1(_02992_),
    .B2(_02999_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _19523_ (.A(_02979_),
    .B(_02989_),
    .X(_03000_));
 sky130_fd_sc_hd__o21ai_1 _19524_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .B1(_02906_),
    .Y(_03001_));
 sky130_fd_sc_hd__xnor2_1 _19525_ (.A(_02906_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_03002_));
 sky130_fd_sc_hd__a21oi_1 _19526_ (.A1(_03000_),
    .A2(_03001_),
    .B1(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__and3_1 _19527_ (.A(_03002_),
    .B(_03000_),
    .C(_03001_),
    .X(_03004_));
 sky130_fd_sc_hd__nor2_1 _19528_ (.A(_03003_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__mux2_1 _19529_ (.A0(_02994_),
    .A1(_02995_),
    .S(_02998_),
    .X(_03006_));
 sky130_fd_sc_hd__or2_1 _19530_ (.A(_04034_),
    .B(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__o221a_1 _19531_ (.A1(\rbzero.wall_tracer.rayAddendY[9] ),
    .A2(_07718_),
    .B1(_07831_),
    .B2(_03005_),
    .C1(_03007_),
    .X(_00819_));
 sky130_fd_sc_hd__nor2_1 _19532_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_02987_),
    .Y(_03008_));
 sky130_fd_sc_hd__or3_1 _19533_ (.A(_02906_),
    .B(_04034_),
    .C(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__a21oi_1 _19534_ (.A1(_02906_),
    .A2(\rbzero.wall_tracer.rayAddendY[9] ),
    .B1(_03003_),
    .Y(_03010_));
 sky130_fd_sc_hd__xnor2_1 _19535_ (.A(_02906_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_03011_));
 sky130_fd_sc_hd__xnor2_1 _19536_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__o2bb2a_1 _19537_ (.A1_N(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2_N(_07695_),
    .B1(_07830_),
    .B2(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__nand2_1 _19538_ (.A(_03009_),
    .B(_03013_),
    .Y(_00820_));
 sky130_fd_sc_hd__or4bb_1 _19539_ (.A(\rbzero.wall_tracer.rayAddendY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .C_N(_03001_),
    .D_N(_02906_),
    .X(_03014_));
 sky130_fd_sc_hd__or3_1 _19540_ (.A(_03002_),
    .B(_03000_),
    .C(_03011_),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _19541_ (.A0(_02906_),
    .A1(_03014_),
    .S(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__nor2_1 _19542_ (.A(_07677_),
    .B(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__xnor2_1 _19543_ (.A(\rbzero.wall_tracer.rayAddendY[11] ),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__o21ai_1 _19544_ (.A1(_03914_),
    .A2(_03018_),
    .B1(_03009_),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2b_2 _19545_ (.A(\rbzero.pov.sclk_buffer[2] ),
    .B_N(\rbzero.pov.sclk_buffer[1] ),
    .Y(_03019_));
 sky130_fd_sc_hd__nor2_2 _19546_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_03555_),
    .Y(_03020_));
 sky130_fd_sc_hd__o21ai_1 _19547_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03019_),
    .B1(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__a21oi_1 _19548_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03019_),
    .B1(_03021_),
    .Y(_00822_));
 sky130_fd_sc_hd__and3_1 _19549_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_03019_),
    .X(_03022_));
 sky130_fd_sc_hd__a21o_1 _19550_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03019_),
    .B1(\rbzero.pov.spi_counter[1] ),
    .X(_03023_));
 sky130_fd_sc_hd__and4bb_1 _19551_ (.A_N(\rbzero.pov.spi_counter[5] ),
    .B_N(\rbzero.pov.spi_counter[4] ),
    .C(\rbzero.pov.spi_counter[3] ),
    .D(\rbzero.pov.spi_counter[6] ),
    .X(_03024_));
 sky130_fd_sc_hd__and4bb_1 _19552_ (.A_N(\rbzero.pov.spi_counter[2] ),
    .B_N(\rbzero.pov.spi_counter[1] ),
    .C(\rbzero.pov.spi_counter[0] ),
    .D(_03024_),
    .X(_03025_));
 sky130_fd_sc_hd__a21boi_1 _19553_ (.A1(_03019_),
    .A2(_03025_),
    .B1_N(_03020_),
    .Y(_03026_));
 sky130_fd_sc_hd__and3b_1 _19554_ (.A_N(_03022_),
    .B(_03023_),
    .C(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _19555_ (.A(_03027_),
    .X(_00823_));
 sky130_fd_sc_hd__and2_1 _19556_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(_03022_),
    .X(_03028_));
 sky130_fd_sc_hd__o21ai_1 _19557_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_03022_),
    .B1(_03020_),
    .Y(_03029_));
 sky130_fd_sc_hd__nor2_1 _19558_ (.A(_03028_),
    .B(_03029_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _19559_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_03028_),
    .Y(_03030_));
 sky130_fd_sc_hd__o211a_1 _19560_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_03028_),
    .B1(_03030_),
    .C1(_03026_),
    .X(_00825_));
 sky130_fd_sc_hd__and3_1 _19561_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_03028_),
    .X(_03031_));
 sky130_fd_sc_hd__a31o_1 _19562_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(\rbzero.pov.spi_counter[2] ),
    .A3(_03022_),
    .B1(\rbzero.pov.spi_counter[4] ),
    .X(_03032_));
 sky130_fd_sc_hd__and3b_1 _19563_ (.A_N(_03031_),
    .B(_03020_),
    .C(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _19564_ (.A(_03033_),
    .X(_00826_));
 sky130_fd_sc_hd__and2_1 _19565_ (.A(\rbzero.pov.spi_counter[5] ),
    .B(_03031_),
    .X(_03034_));
 sky130_fd_sc_hd__o21ai_1 _19566_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_03031_),
    .B1(_03020_),
    .Y(_03035_));
 sky130_fd_sc_hd__nor2_1 _19567_ (.A(_03034_),
    .B(_03035_),
    .Y(_00827_));
 sky130_fd_sc_hd__a21boi_1 _19568_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03034_),
    .B1_N(_03026_),
    .Y(_03036_));
 sky130_fd_sc_hd__o21a_1 _19569_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03034_),
    .B1(_03036_),
    .X(_00828_));
 sky130_fd_sc_hd__buf_1 _19570_ (.A(clknet_1_0__leaf__04835_),
    .X(_03037_));
 sky130_fd_sc_hd__buf_1 _19571_ (.A(clknet_1_0__leaf__03037_),
    .X(_03038_));
 sky130_fd_sc_hd__inv_2 _19573__30 (.A(clknet_1_1__leaf__03038_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _19574__31 (.A(clknet_1_1__leaf__03038_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _19575__32 (.A(clknet_1_1__leaf__03038_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _19576__33 (.A(clknet_1_1__leaf__03038_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _19577__34 (.A(clknet_1_0__leaf__03038_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _19578__35 (.A(clknet_1_0__leaf__03038_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _19579__36 (.A(clknet_1_0__leaf__03038_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _19580__37 (.A(clknet_1_0__leaf__03038_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _19581__38 (.A(clknet_1_0__leaf__03038_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _19583__39 (.A(clknet_1_1__leaf__03039_),
    .Y(net160));
 sky130_fd_sc_hd__buf_1 _19582_ (.A(clknet_1_0__leaf__03037_),
    .X(_03039_));
 sky130_fd_sc_hd__inv_2 _19584__40 (.A(clknet_1_1__leaf__03039_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _19585__41 (.A(clknet_1_1__leaf__03039_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _19586__42 (.A(clknet_1_1__leaf__03039_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _19587__43 (.A(clknet_1_1__leaf__03039_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _19588__44 (.A(clknet_1_0__leaf__03039_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _19589__45 (.A(clknet_1_0__leaf__03039_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _19590__46 (.A(clknet_1_0__leaf__03039_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _19591__47 (.A(clknet_1_0__leaf__03039_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _19592__48 (.A(clknet_1_0__leaf__03039_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _19594__49 (.A(clknet_1_1__leaf__03040_),
    .Y(net170));
 sky130_fd_sc_hd__buf_1 _19593_ (.A(clknet_1_0__leaf__03037_),
    .X(_03040_));
 sky130_fd_sc_hd__inv_2 _19595__50 (.A(clknet_1_1__leaf__03040_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _19596__51 (.A(clknet_1_0__leaf__03040_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _19597__52 (.A(clknet_1_0__leaf__03040_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _19598__53 (.A(clknet_1_0__leaf__03040_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _19599__54 (.A(clknet_1_0__leaf__03040_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _19600__55 (.A(clknet_1_0__leaf__03040_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _19601__56 (.A(clknet_1_0__leaf__03040_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _19602__57 (.A(clknet_1_1__leaf__03040_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _19603__58 (.A(clknet_1_1__leaf__03040_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _19605__59 (.A(clknet_1_0__leaf__03041_),
    .Y(net180));
 sky130_fd_sc_hd__buf_1 _19604_ (.A(clknet_1_0__leaf__03037_),
    .X(_03041_));
 sky130_fd_sc_hd__inv_2 _19606__60 (.A(clknet_1_0__leaf__03041_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _19607__61 (.A(clknet_1_1__leaf__03041_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _19608__62 (.A(clknet_1_1__leaf__03041_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _19609__63 (.A(clknet_1_1__leaf__03041_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _19610__64 (.A(clknet_1_1__leaf__03041_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _19611__65 (.A(clknet_1_0__leaf__03041_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _19612__66 (.A(clknet_1_0__leaf__03041_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _19613__67 (.A(clknet_1_0__leaf__03041_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _19614__68 (.A(clknet_1_0__leaf__03041_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _19616__69 (.A(clknet_1_0__leaf__03042_),
    .Y(net190));
 sky130_fd_sc_hd__buf_1 _19615_ (.A(clknet_1_1__leaf__03037_),
    .X(_03042_));
 sky130_fd_sc_hd__inv_2 _19617__70 (.A(clknet_1_0__leaf__03042_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _19618__71 (.A(clknet_1_0__leaf__03042_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _19619__72 (.A(clknet_1_0__leaf__03042_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _19620__73 (.A(clknet_1_1__leaf__03042_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _19621__74 (.A(clknet_1_1__leaf__03042_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _19622__75 (.A(clknet_1_1__leaf__03042_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _19623__76 (.A(clknet_1_1__leaf__03042_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _19624__77 (.A(clknet_1_0__leaf__03042_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _19625__78 (.A(clknet_1_1__leaf__03042_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _19627__79 (.A(clknet_1_0__leaf__03043_),
    .Y(net200));
 sky130_fd_sc_hd__buf_1 _19626_ (.A(clknet_1_1__leaf__03037_),
    .X(_03043_));
 sky130_fd_sc_hd__inv_2 _19628__80 (.A(clknet_1_0__leaf__03043_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _19629__81 (.A(clknet_1_1__leaf__03043_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _19630__82 (.A(clknet_1_1__leaf__03043_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _19631__83 (.A(clknet_1_1__leaf__03043_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _19632__84 (.A(clknet_1_1__leaf__03043_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _19633__85 (.A(clknet_1_1__leaf__03043_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _19634__86 (.A(clknet_1_1__leaf__03043_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _19635__87 (.A(clknet_1_0__leaf__03043_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _19636__88 (.A(clknet_1_0__leaf__03043_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _19639__89 (.A(clknet_1_0__leaf__03045_),
    .Y(net210));
 sky130_fd_sc_hd__buf_1 _19637_ (.A(clknet_1_0__leaf__04835_),
    .X(_03044_));
 sky130_fd_sc_hd__buf_1 _19638_ (.A(clknet_1_1__leaf__03044_),
    .X(_03045_));
 sky130_fd_sc_hd__inv_2 _19640__90 (.A(clknet_1_0__leaf__03045_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _19641__91 (.A(clknet_1_0__leaf__03045_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _19642__92 (.A(clknet_1_1__leaf__03045_),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _20055__93 (.A(clknet_1_1__leaf__03045_),
    .Y(net214));
 sky130_fd_sc_hd__nand2_1 _19643_ (.A(_03020_),
    .B(_03019_),
    .Y(_03046_));
 sky130_fd_sc_hd__buf_4 _19644_ (.A(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_4 _19645_ (.A(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _19646_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _19647_ (.A(_03049_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _19648_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_03048_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _19649_ (.A(_03050_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _19650_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_03048_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _19651_ (.A(_03051_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _19652_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_03048_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _19653_ (.A(_03052_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _19654_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_03048_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _19655_ (.A(_03053_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _19656_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_03048_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _19657_ (.A(_03054_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _19658_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_03048_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _19659_ (.A(_03055_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _19660_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_03048_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _19661_ (.A(_03056_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _19662_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_03048_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _19663_ (.A(_03057_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _19664_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_03048_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _19665_ (.A(_03058_),
    .X(_00902_));
 sky130_fd_sc_hd__clkbuf_4 _19666_ (.A(_03047_),
    .X(_03059_));
 sky130_fd_sc_hd__mux2_1 _19667_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _19668_ (.A(_03060_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _19669_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_03059_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _19670_ (.A(_03061_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19671_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_03059_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _19672_ (.A(_03062_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _19673_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_03059_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _19674_ (.A(_03063_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19675_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_03059_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _19676_ (.A(_03064_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19677_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_03059_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _19678_ (.A(_03065_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _19679_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_03059_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _19680_ (.A(_03066_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _19681_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_03059_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _19682_ (.A(_03067_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _19683_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_03059_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _19684_ (.A(_03068_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19685_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_03059_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _19686_ (.A(_03069_),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_4 _19687_ (.A(_03047_),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _19688_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_1 _19689_ (.A(_03071_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _19690_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_03070_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _19691_ (.A(_03072_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _19692_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_03070_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _19693_ (.A(_03073_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _19694_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_03070_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _19695_ (.A(_03074_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _19696_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_03070_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _19697_ (.A(_03075_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _19698_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_03070_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _19699_ (.A(_03076_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _19700_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_03070_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_1 _19701_ (.A(_03077_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _19702_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_03070_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _19703_ (.A(_03078_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _19704_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_03070_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _19705_ (.A(_03079_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _19706_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_03070_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _19707_ (.A(_03080_),
    .X(_00922_));
 sky130_fd_sc_hd__buf_4 _19708_ (.A(_03047_),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _19709_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _19710_ (.A(_03082_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _19711_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_03081_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _19712_ (.A(_03083_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _19713_ (.A0(net512),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_03081_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_1 _19714_ (.A(_03084_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _19715_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_03081_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _19716_ (.A(_03085_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _19717_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_03081_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _19718_ (.A(_03086_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19719_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_03081_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _19720_ (.A(_03087_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _19721_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_03081_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _19722_ (.A(_03088_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19723_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_03081_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_1 _19724_ (.A(_03089_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19725_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_03081_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _19726_ (.A(_03090_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _19727_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_03081_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _19728_ (.A(_03091_),
    .X(_00932_));
 sky130_fd_sc_hd__clkbuf_4 _19729_ (.A(_03047_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _19730_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _19731_ (.A(_03093_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _19732_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_03092_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_1 _19733_ (.A(_03094_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _19734_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_03092_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_1 _19735_ (.A(_03095_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _19736_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_03092_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _19737_ (.A(_03096_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19738_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_03092_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _19739_ (.A(_03097_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _19740_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_03092_),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _19741_ (.A(_03098_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _19742_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_03092_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _19743_ (.A(_03099_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19744_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_03092_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _19745_ (.A(_03100_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19746_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_03092_),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _19747_ (.A(_03101_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _19748_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_03092_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _19749_ (.A(_03102_),
    .X(_00942_));
 sky130_fd_sc_hd__clkbuf_4 _19750_ (.A(_03047_),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _19751_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _19752_ (.A(_03104_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _19753_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_03103_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _19754_ (.A(_03105_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _19755_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_03103_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _19756_ (.A(_03106_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _19757_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_03103_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _19758_ (.A(_03107_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _19759_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_03103_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _19760_ (.A(_03108_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _19761_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_03103_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _19762_ (.A(_03109_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _19763_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_03103_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _19764_ (.A(_03110_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _19765_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_03103_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _19766_ (.A(_03111_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _19767_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_03103_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _19768_ (.A(_03112_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _19769_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_03103_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_1 _19770_ (.A(_03113_),
    .X(_00952_));
 sky130_fd_sc_hd__buf_4 _19771_ (.A(_03046_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _19772_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _19773_ (.A(_03115_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _19774_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_03114_),
    .X(_03116_));
 sky130_fd_sc_hd__clkbuf_1 _19775_ (.A(_03116_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _19776_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_03114_),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_1 _19777_ (.A(_03117_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _19778_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_03114_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _19779_ (.A(_03118_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _19780_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_03114_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _19781_ (.A(_03119_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19782_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_03114_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _19783_ (.A(_03120_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19784_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_03114_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _19785_ (.A(_03121_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19786_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_03114_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_1 _19787_ (.A(_03122_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _19788_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_03114_),
    .X(_03123_));
 sky130_fd_sc_hd__clkbuf_1 _19789_ (.A(_03123_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _19790_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_03114_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _19791_ (.A(_03124_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _19792_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_03047_),
    .X(_03125_));
 sky130_fd_sc_hd__clkbuf_1 _19793_ (.A(_03125_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _19794_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_03047_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _19795_ (.A(_03126_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _19796_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_03047_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _19797_ (.A(_03127_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _19798_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_03047_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _19799_ (.A(_03128_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _19800_ (.A0(_04867_),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_02695_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _19801_ (.A(_03129_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _19802_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_05189_),
    .X(_03130_));
 sky130_fd_sc_hd__clkbuf_1 _19803_ (.A(_03130_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _19804_ (.A0(net50),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_02695_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_1 _19805_ (.A(_03131_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _19806_ (.A0(\rbzero.pov.ss_buffer[1] ),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_05189_),
    .X(_03132_));
 sky130_fd_sc_hd__clkbuf_1 _19807_ (.A(_03132_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _19808_ (.A0(net52),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_02695_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_1 _19809_ (.A(_03133_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _19810_ (.A0(\rbzero.pov.sclk_buffer[1] ),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_05189_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_1 _19811_ (.A(_03134_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19812_ (.A0(\rbzero.pov.sclk_buffer[2] ),
    .A1(\rbzero.pov.sclk_buffer[1] ),
    .S(_05189_),
    .X(_03135_));
 sky130_fd_sc_hd__clkbuf_1 _19813_ (.A(_03135_),
    .X(_00973_));
 sky130_fd_sc_hd__and2_1 _19814_ (.A(\rbzero.pov.ready ),
    .B(_02821_),
    .X(_03136_));
 sky130_fd_sc_hd__buf_2 _19815_ (.A(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__o21ai_2 _19816_ (.A1(net38),
    .A2(_03137_),
    .B1(_02708_),
    .Y(_03138_));
 sky130_fd_sc_hd__clkbuf_4 _19817_ (.A(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__inv_2 _19818_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_03140_));
 sky130_fd_sc_hd__clkbuf_4 _19819_ (.A(_02822_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_1 _19820_ (.A0(_03140_),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_4 _19821_ (.A(_03138_),
    .X(_03143_));
 sky130_fd_sc_hd__nand2_1 _19822_ (.A(_03140_),
    .B(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__o211a_1 _19823_ (.A1(_03139_),
    .A2(_03142_),
    .B1(_03144_),
    .C1(_02765_),
    .X(_00974_));
 sky130_fd_sc_hd__nor2_1 _19824_ (.A(_02728_),
    .B(_02820_),
    .Y(_03145_));
 sky130_fd_sc_hd__buf_4 _19825_ (.A(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _19826_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(_07985_),
    .S(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__inv_2 _19827_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_1 _19828_ (.A(_03148_),
    .B(_03143_),
    .Y(_03149_));
 sky130_fd_sc_hd__o211a_1 _19829_ (.A1(_03139_),
    .A2(_03147_),
    .B1(_03149_),
    .C1(_02765_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _19830_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(_07999_),
    .S(_03146_),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _19831_ (.A(_08000_),
    .B(_03143_),
    .Y(_03151_));
 sky130_fd_sc_hd__o211a_1 _19832_ (.A1(_03139_),
    .A2(_03150_),
    .B1(_03151_),
    .C1(_02765_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _19833_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(_07900_),
    .S(_03146_),
    .X(_03152_));
 sky130_fd_sc_hd__nand2_1 _19834_ (.A(_07901_),
    .B(_03143_),
    .Y(_03153_));
 sky130_fd_sc_hd__o211a_1 _19835_ (.A1(_03139_),
    .A2(_03152_),
    .B1(_03153_),
    .C1(_02765_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _19836_ (.A0(\rbzero.pov.ready_buffer[63] ),
    .A1(_07914_),
    .S(_03146_),
    .X(_03154_));
 sky130_fd_sc_hd__o21a_2 _19837_ (.A1(net38),
    .A2(_03137_),
    .B1(_02708_),
    .X(_03155_));
 sky130_fd_sc_hd__or2_1 _19838_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_4 _19839_ (.A(_05190_),
    .X(_03157_));
 sky130_fd_sc_hd__o211a_1 _19840_ (.A1(_03139_),
    .A2(_03154_),
    .B1(_03156_),
    .C1(_03157_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _19841_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_07948_),
    .S(_03146_),
    .X(_03158_));
 sky130_fd_sc_hd__nand2_1 _19842_ (.A(_07949_),
    .B(_03143_),
    .Y(_03159_));
 sky130_fd_sc_hd__o211a_1 _19843_ (.A1(_03139_),
    .A2(_03158_),
    .B1(_03159_),
    .C1(_03157_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _19844_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(_08066_),
    .S(_03146_),
    .X(_03160_));
 sky130_fd_sc_hd__nand2_1 _19845_ (.A(_08067_),
    .B(_03143_),
    .Y(_03161_));
 sky130_fd_sc_hd__o211a_1 _19846_ (.A1(_03139_),
    .A2(_03160_),
    .B1(_03161_),
    .C1(_03157_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _19847_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(_08077_),
    .S(_03146_),
    .X(_03162_));
 sky130_fd_sc_hd__nand2_1 _19848_ (.A(_08078_),
    .B(_03143_),
    .Y(_03163_));
 sky130_fd_sc_hd__o211a_1 _19849_ (.A1(_03139_),
    .A2(_03162_),
    .B1(_03163_),
    .C1(_03157_),
    .X(_00981_));
 sky130_fd_sc_hd__clkbuf_4 _19850_ (.A(_03146_),
    .X(_03164_));
 sky130_fd_sc_hd__nor2_1 _19851_ (.A(\rbzero.pov.ready_buffer[67] ),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__a211oi_1 _19852_ (.A1(_08093_),
    .A2(_03164_),
    .B1(_03143_),
    .C1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__a211o_1 _19853_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_03139_),
    .B1(_03166_),
    .C1(net60),
    .X(_00982_));
 sky130_fd_sc_hd__or2_1 _19854_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08028_),
    .X(_03167_));
 sky130_fd_sc_hd__nand2_1 _19855_ (.A(_03145_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__a21o_1 _19856_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_08028_),
    .B1(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__o211a_1 _19857_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_03164_),
    .B1(_03155_),
    .C1(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__a211o_1 _19858_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03139_),
    .B1(_03170_),
    .C1(net60),
    .X(_00983_));
 sky130_fd_sc_hd__nor2_1 _19859_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03167_),
    .Y(_03171_));
 sky130_fd_sc_hd__and2_1 _19860_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03167_),
    .X(_03172_));
 sky130_fd_sc_hd__or2_1 _19861_ (.A(\rbzero.pov.ready_buffer[69] ),
    .B(_03145_),
    .X(_03173_));
 sky130_fd_sc_hd__o311a_1 _19862_ (.A1(_03141_),
    .A2(_03171_),
    .A3(_03172_),
    .B1(_03173_),
    .C1(_03155_),
    .X(_03174_));
 sky130_fd_sc_hd__buf_4 _19863_ (.A(_03911_),
    .X(_03175_));
 sky130_fd_sc_hd__a211o_1 _19864_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03143_),
    .B1(_03174_),
    .C1(_03175_),
    .X(_00984_));
 sky130_fd_sc_hd__or3_1 _19865_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(\rbzero.debug_overlay.playerX[1] ),
    .C(_03167_),
    .X(_03176_));
 sky130_fd_sc_hd__o21ai_1 _19866_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03167_),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .Y(_03177_));
 sky130_fd_sc_hd__a21oi_1 _19867_ (.A1(_03176_),
    .A2(_03177_),
    .B1(_02822_),
    .Y(_03178_));
 sky130_fd_sc_hd__a211o_1 _19868_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_02823_),
    .B1(_03138_),
    .C1(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__o211a_1 _19869_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03155_),
    .B1(_03179_),
    .C1(_03157_),
    .X(_00985_));
 sky130_fd_sc_hd__nor2_1 _19870_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03176_),
    .Y(_03180_));
 sky130_fd_sc_hd__a21o_1 _19871_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03176_),
    .B1(_02822_),
    .X(_03181_));
 sky130_fd_sc_hd__o221a_1 _19872_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_03146_),
    .B1(_03180_),
    .B2(_03181_),
    .C1(_03155_),
    .X(_03182_));
 sky130_fd_sc_hd__a211o_1 _19873_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03143_),
    .B1(_03182_),
    .C1(_03175_),
    .X(_00986_));
 sky130_fd_sc_hd__nor2_1 _19874_ (.A(_02820_),
    .B(_03180_),
    .Y(_03183_));
 sky130_fd_sc_hd__o21a_1 _19875_ (.A1(_03138_),
    .A2(_03183_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .X(_03184_));
 sky130_fd_sc_hd__and2b_1 _19876_ (.A_N(\rbzero.debug_overlay.playerX[4] ),
    .B(_03180_),
    .X(_03185_));
 sky130_fd_sc_hd__o21a_1 _19877_ (.A1(_02820_),
    .A2(_03185_),
    .B1(_03155_),
    .X(_03186_));
 sky130_fd_sc_hd__o21a_1 _19878_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_03164_),
    .B1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__o21a_1 _19879_ (.A1(_03184_),
    .A2(_03187_),
    .B1(_02714_),
    .X(_00987_));
 sky130_fd_sc_hd__inv_2 _19880_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .Y(_03188_));
 sky130_fd_sc_hd__nor2_1 _19881_ (.A(_03188_),
    .B(_03186_),
    .Y(_03189_));
 sky130_fd_sc_hd__a21o_1 _19882_ (.A1(_03188_),
    .A2(_03185_),
    .B1(_02822_),
    .X(_03190_));
 sky130_fd_sc_hd__o211a_1 _19883_ (.A1(\rbzero.pov.ready_buffer[73] ),
    .A2(_03164_),
    .B1(_03155_),
    .C1(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__o21a_1 _19884_ (.A1(_03189_),
    .A2(_03191_),
    .B1(_02714_),
    .X(_00988_));
 sky130_fd_sc_hd__o21ai_2 _19885_ (.A1(net39),
    .A2(_03137_),
    .B1(_02708_),
    .Y(_03192_));
 sky130_fd_sc_hd__clkbuf_4 _19886_ (.A(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__inv_2 _19887_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_03194_));
 sky130_fd_sc_hd__mux2_1 _19888_ (.A0(_03194_),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_02822_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2_1 _19889_ (.A(_03194_),
    .B(_03193_),
    .Y(_03196_));
 sky130_fd_sc_hd__o211a_1 _19890_ (.A1(_03193_),
    .A2(_03195_),
    .B1(_03196_),
    .C1(_03157_),
    .X(_00989_));
 sky130_fd_sc_hd__o21a_1 _19891_ (.A1(net39),
    .A2(_03137_),
    .B1(_02708_),
    .X(_03197_));
 sky130_fd_sc_hd__buf_2 _19892_ (.A(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__nand2_1 _19893_ (.A(\rbzero.pov.ready_buffer[45] ),
    .B(_02823_),
    .Y(_03199_));
 sky130_fd_sc_hd__o211ai_1 _19894_ (.A1(_07982_),
    .A2(_02823_),
    .B1(_03198_),
    .C1(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o211a_1 _19895_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(_03198_),
    .B1(_03200_),
    .C1(_03157_),
    .X(_00990_));
 sky130_fd_sc_hd__nor2_1 _19896_ (.A(_08004_),
    .B(_03141_),
    .Y(_03201_));
 sky130_fd_sc_hd__a211o_1 _19897_ (.A1(\rbzero.pov.ready_buffer[46] ),
    .A2(_02823_),
    .B1(_03193_),
    .C1(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__o211a_1 _19898_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_03198_),
    .B1(_03202_),
    .C1(_03157_),
    .X(_00991_));
 sky130_fd_sc_hd__nor2_1 _19899_ (.A(_07908_),
    .B(_03141_),
    .Y(_03203_));
 sky130_fd_sc_hd__a211o_1 _19900_ (.A1(\rbzero.pov.ready_buffer[47] ),
    .A2(_02823_),
    .B1(_03193_),
    .C1(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__o211a_1 _19901_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_03198_),
    .B1(_03204_),
    .C1(_03157_),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_1 _19902_ (.A(_07917_),
    .B(_03141_),
    .Y(_03205_));
 sky130_fd_sc_hd__a211o_1 _19903_ (.A1(\rbzero.pov.ready_buffer[48] ),
    .A2(_02823_),
    .B1(_03193_),
    .C1(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__o211a_1 _19904_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_03198_),
    .B1(_03206_),
    .C1(_03157_),
    .X(_00993_));
 sky130_fd_sc_hd__nor2_1 _19905_ (.A(_07954_),
    .B(_03141_),
    .Y(_03207_));
 sky130_fd_sc_hd__a211o_1 _19906_ (.A1(\rbzero.pov.ready_buffer[49] ),
    .A2(_02823_),
    .B1(_03192_),
    .C1(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__buf_6 _19907_ (.A(_05190_),
    .X(_03209_));
 sky130_fd_sc_hd__o211a_1 _19908_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_03198_),
    .B1(_03208_),
    .C1(_03209_),
    .X(_00994_));
 sky130_fd_sc_hd__nor2_1 _19909_ (.A(_08070_),
    .B(_03141_),
    .Y(_03210_));
 sky130_fd_sc_hd__a211o_1 _19910_ (.A1(\rbzero.pov.ready_buffer[50] ),
    .A2(_03141_),
    .B1(_03192_),
    .C1(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__o211a_1 _19911_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_03198_),
    .B1(_03211_),
    .C1(_03209_),
    .X(_00995_));
 sky130_fd_sc_hd__nand2_1 _19912_ (.A(\rbzero.pov.ready_buffer[51] ),
    .B(_02823_),
    .Y(_03212_));
 sky130_fd_sc_hd__o211ai_1 _19913_ (.A1(_08080_),
    .A2(_02823_),
    .B1(_03197_),
    .C1(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__o211a_1 _19914_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_03198_),
    .B1(_03213_),
    .C1(_03209_),
    .X(_00996_));
 sky130_fd_sc_hd__nor2_1 _19915_ (.A(\rbzero.pov.ready_buffer[52] ),
    .B(_03164_),
    .Y(_03214_));
 sky130_fd_sc_hd__a211oi_1 _19916_ (.A1(_08089_),
    .A2(_03164_),
    .B1(_03193_),
    .C1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__a211o_1 _19917_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_03193_),
    .B1(_03215_),
    .C1(_03175_),
    .X(_00997_));
 sky130_fd_sc_hd__or2_1 _19918_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08030_),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_1 _19919_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08030_),
    .Y(_03217_));
 sky130_fd_sc_hd__a21oi_1 _19920_ (.A1(_03216_),
    .A2(_03217_),
    .B1(_02822_),
    .Y(_03218_));
 sky130_fd_sc_hd__a211o_1 _19921_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_03141_),
    .B1(_03192_),
    .C1(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__o211a_1 _19922_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03198_),
    .B1(_03219_),
    .C1(_03209_),
    .X(_00998_));
 sky130_fd_sc_hd__o21ai_1 _19923_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03216_),
    .B1(_03145_),
    .Y(_03220_));
 sky130_fd_sc_hd__a21o_1 _19924_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03216_),
    .B1(_03220_),
    .X(_03221_));
 sky130_fd_sc_hd__o211a_1 _19925_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_03164_),
    .B1(_03197_),
    .C1(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__a211o_1 _19926_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03193_),
    .B1(_03222_),
    .C1(_03175_),
    .X(_00999_));
 sky130_fd_sc_hd__or3_1 _19927_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .C(_03216_),
    .X(_03223_));
 sky130_fd_sc_hd__o21ai_1 _19928_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03216_),
    .B1(\rbzero.debug_overlay.playerY[2] ),
    .Y(_03224_));
 sky130_fd_sc_hd__a21oi_1 _19929_ (.A1(_03223_),
    .A2(_03224_),
    .B1(_02822_),
    .Y(_03225_));
 sky130_fd_sc_hd__a211o_1 _19930_ (.A1(\rbzero.pov.ready_buffer[55] ),
    .A2(_03141_),
    .B1(_03192_),
    .C1(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__o211a_1 _19931_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_03198_),
    .B1(_03226_),
    .C1(_03209_),
    .X(_01000_));
 sky130_fd_sc_hd__nor2_1 _19932_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .B(_03223_),
    .Y(_03227_));
 sky130_fd_sc_hd__a21o_1 _19933_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03223_),
    .B1(_02822_),
    .X(_03228_));
 sky130_fd_sc_hd__o221a_1 _19934_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_03146_),
    .B1(_03227_),
    .B2(_03228_),
    .C1(_03197_),
    .X(_03229_));
 sky130_fd_sc_hd__a211o_1 _19935_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03193_),
    .B1(_03229_),
    .C1(_03175_),
    .X(_01001_));
 sky130_fd_sc_hd__nor2_1 _19936_ (.A(_02820_),
    .B(_03227_),
    .Y(_03230_));
 sky130_fd_sc_hd__o21a_1 _19937_ (.A1(_03193_),
    .A2(_03230_),
    .B1(\rbzero.debug_overlay.playerY[4] ),
    .X(_03231_));
 sky130_fd_sc_hd__and2_1 _19938_ (.A(_03920_),
    .B(_03227_),
    .X(_03232_));
 sky130_fd_sc_hd__o21a_1 _19939_ (.A1(_02820_),
    .A2(_03232_),
    .B1(_03197_),
    .X(_03233_));
 sky130_fd_sc_hd__o21a_1 _19940_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_03164_),
    .B1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__o21a_1 _19941_ (.A1(_03231_),
    .A2(_03234_),
    .B1(_02714_),
    .X(_01002_));
 sky130_fd_sc_hd__inv_2 _19942_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .Y(_03235_));
 sky130_fd_sc_hd__nor2_1 _19943_ (.A(_03235_),
    .B(_03233_),
    .Y(_03236_));
 sky130_fd_sc_hd__a31o_1 _19944_ (.A1(_03235_),
    .A2(_03920_),
    .A3(_03227_),
    .B1(_02822_),
    .X(_03237_));
 sky130_fd_sc_hd__o211a_1 _19945_ (.A1(\rbzero.pov.ready_buffer[58] ),
    .A2(_03164_),
    .B1(_03197_),
    .C1(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__o21a_1 _19946_ (.A1(_03236_),
    .A2(_03238_),
    .B1(_02714_),
    .X(_01003_));
 sky130_fd_sc_hd__nand3_4 _19947_ (.A(\rbzero.pov.ready ),
    .B(_02708_),
    .C(_02820_),
    .Y(_03239_));
 sky130_fd_sc_hd__buf_2 _19948_ (.A(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__and3_1 _19949_ (.A(\rbzero.pov.ready ),
    .B(_02707_),
    .C(_02820_),
    .X(_03241_));
 sky130_fd_sc_hd__buf_2 _19950_ (.A(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__buf_2 _19951_ (.A(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__o221a_1 _19952_ (.A1(\rbzero.pov.ready_buffer[33] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .C1(_03209_),
    .X(_01004_));
 sky130_fd_sc_hd__o221a_1 _19953_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[-8] ),
    .C1(_03209_),
    .X(_01005_));
 sky130_fd_sc_hd__o221a_1 _19954_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .C1(_03209_),
    .X(_01006_));
 sky130_fd_sc_hd__buf_2 _19955_ (.A(_02721_),
    .X(_03244_));
 sky130_fd_sc_hd__o221a_1 _19956_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[-6] ),
    .C1(_03244_),
    .X(_01007_));
 sky130_fd_sc_hd__and3_1 _19957_ (.A(\rbzero.pov.ready ),
    .B(_02707_),
    .C(_02820_),
    .X(_03245_));
 sky130_fd_sc_hd__clkbuf_4 _19958_ (.A(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_4 _19959_ (.A(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__nand2_4 _19960_ (.A(_02708_),
    .B(_03137_),
    .Y(_03248_));
 sky130_fd_sc_hd__clkbuf_4 _19961_ (.A(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_6 _19962_ (.A(_02695_),
    .X(_03250_));
 sky130_fd_sc_hd__a221o_1 _19963_ (.A1(\rbzero.pov.ready_buffer[37] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingX[-5] ),
    .C1(_03250_),
    .X(_01008_));
 sky130_fd_sc_hd__a221o_1 _19964_ (.A1(\rbzero.pov.ready_buffer[38] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingX[-4] ),
    .C1(_03250_),
    .X(_01009_));
 sky130_fd_sc_hd__clkbuf_4 _19965_ (.A(_02695_),
    .X(_03251_));
 sky130_fd_sc_hd__a221o_1 _19966_ (.A1(\rbzero.pov.ready_buffer[39] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingX[-3] ),
    .C1(_03251_),
    .X(_01010_));
 sky130_fd_sc_hd__o221a_1 _19967_ (.A1(\rbzero.pov.ready_buffer[40] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[-2] ),
    .C1(_03244_),
    .X(_01011_));
 sky130_fd_sc_hd__a221o_1 _19968_ (.A1(\rbzero.pov.ready_buffer[41] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingX[-1] ),
    .C1(_03251_),
    .X(_01012_));
 sky130_fd_sc_hd__o221a_1 _19969_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .C1(_03244_),
    .X(_01013_));
 sky130_fd_sc_hd__o221a_1 _19970_ (.A1(\rbzero.pov.ready_buffer[43] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingX[10] ),
    .C1(_03244_),
    .X(_01014_));
 sky130_fd_sc_hd__o221a_1 _19971_ (.A1(\rbzero.pov.ready_buffer[22] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .C1(_03244_),
    .X(_01015_));
 sky130_fd_sc_hd__o221a_1 _19972_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingY[-8] ),
    .C1(_03244_),
    .X(_01016_));
 sky130_fd_sc_hd__a221o_1 _19973_ (.A1(\rbzero.pov.ready_buffer[24] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .C1(_03251_),
    .X(_01017_));
 sky130_fd_sc_hd__a221o_1 _19974_ (.A1(\rbzero.pov.ready_buffer[25] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingY[-6] ),
    .C1(_03251_),
    .X(_01018_));
 sky130_fd_sc_hd__a221o_1 _19975_ (.A1(\rbzero.pov.ready_buffer[26] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .C1(_03251_),
    .X(_01019_));
 sky130_fd_sc_hd__o221a_1 _19976_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_03240_),
    .B1(_03243_),
    .B2(\rbzero.debug_overlay.facingY[-4] ),
    .C1(_03244_),
    .X(_01020_));
 sky130_fd_sc_hd__clkbuf_4 _19977_ (.A(_03239_),
    .X(_03252_));
 sky130_fd_sc_hd__buf_2 _19978_ (.A(_03242_),
    .X(_03253_));
 sky130_fd_sc_hd__o221a_1 _19979_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .C1(_03244_),
    .X(_01021_));
 sky130_fd_sc_hd__a221o_1 _19980_ (.A1(net513),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .C1(_03251_),
    .X(_01022_));
 sky130_fd_sc_hd__o221a_1 _19981_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .C1(_03244_),
    .X(_01023_));
 sky130_fd_sc_hd__a221o_1 _19982_ (.A1(net70),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingY[0] ),
    .C1(_03251_),
    .X(_01024_));
 sky130_fd_sc_hd__a221o_1 _19983_ (.A1(\rbzero.pov.ready_buffer[32] ),
    .A2(_03247_),
    .B1(_03249_),
    .B2(\rbzero.debug_overlay.facingY[10] ),
    .C1(_03251_),
    .X(_01025_));
 sky130_fd_sc_hd__a221o_1 _19984_ (.A1(\rbzero.pov.ready_buffer[11] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneX[-9] ),
    .C1(_03251_),
    .X(_01026_));
 sky130_fd_sc_hd__o221a_1 _19985_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(\rbzero.debug_overlay.vplaneX[-8] ),
    .C1(_03244_),
    .X(_01027_));
 sky130_fd_sc_hd__clkbuf_4 _19986_ (.A(_02721_),
    .X(_03254_));
 sky130_fd_sc_hd__o221a_1 _19987_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .C1(_03254_),
    .X(_01028_));
 sky130_fd_sc_hd__o221a_1 _19988_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(\rbzero.debug_overlay.vplaneX[-6] ),
    .C1(_03254_),
    .X(_01029_));
 sky130_fd_sc_hd__a221o_1 _19989_ (.A1(\rbzero.pov.ready_buffer[15] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneX[-5] ),
    .C1(_03251_),
    .X(_01030_));
 sky130_fd_sc_hd__a221o_1 _19990_ (.A1(\rbzero.pov.ready_buffer[16] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneX[-4] ),
    .C1(_02741_),
    .X(_01031_));
 sky130_fd_sc_hd__o221a_1 _19991_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(_04462_),
    .C1(_03254_),
    .X(_01032_));
 sky130_fd_sc_hd__a221o_1 _19992_ (.A1(\rbzero.pov.ready_buffer[18] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .C1(_02741_),
    .X(_01033_));
 sky130_fd_sc_hd__o221a_1 _19993_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(_07730_),
    .C1(_03254_),
    .X(_01034_));
 sky130_fd_sc_hd__o221a_1 _19994_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(_07742_),
    .C1(_03254_),
    .X(_01035_));
 sky130_fd_sc_hd__o221a_1 _19995_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(_07821_),
    .C1(_03254_),
    .X(_01036_));
 sky130_fd_sc_hd__o221a_1 _19996_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_03252_),
    .B1(_03253_),
    .B2(\rbzero.debug_overlay.vplaneY[-9] ),
    .C1(_03254_),
    .X(_01037_));
 sky130_fd_sc_hd__o221a_1 _19997_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_03239_),
    .B1(_03242_),
    .B2(\rbzero.debug_overlay.vplaneY[-8] ),
    .C1(_03254_),
    .X(_01038_));
 sky130_fd_sc_hd__o221a_1 _19998_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_03239_),
    .B1(_03242_),
    .B2(\rbzero.debug_overlay.vplaneY[-7] ),
    .C1(_03254_),
    .X(_01039_));
 sky130_fd_sc_hd__a221o_1 _19999_ (.A1(\rbzero.pov.ready_buffer[3] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneY[-6] ),
    .C1(_02741_),
    .X(_01040_));
 sky130_fd_sc_hd__a221o_1 _20000_ (.A1(\rbzero.pov.ready_buffer[4] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneY[-5] ),
    .C1(_02741_),
    .X(_01041_));
 sky130_fd_sc_hd__a221o_1 _20001_ (.A1(\rbzero.pov.ready_buffer[5] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneY[-4] ),
    .C1(_02741_),
    .X(_01042_));
 sky130_fd_sc_hd__o221a_1 _20002_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_03239_),
    .B1(_03242_),
    .B2(_04471_),
    .C1(_03254_),
    .X(_01043_));
 sky130_fd_sc_hd__a221o_1 _20003_ (.A1(\rbzero.pov.ready_buffer[7] ),
    .A2(_03246_),
    .B1(_03248_),
    .B2(\rbzero.debug_overlay.vplaneY[-2] ),
    .C1(_02741_),
    .X(_01044_));
 sky130_fd_sc_hd__o221a_1 _20004_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_03239_),
    .B1(_03242_),
    .B2(\rbzero.debug_overlay.vplaneY[-1] ),
    .C1(_02730_),
    .X(_01045_));
 sky130_fd_sc_hd__o221a_1 _20005_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_03239_),
    .B1(_03242_),
    .B2(\rbzero.debug_overlay.vplaneY[0] ),
    .C1(_02730_),
    .X(_01046_));
 sky130_fd_sc_hd__o221a_1 _20006_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_03239_),
    .B1(_03242_),
    .B2(_02906_),
    .C1(_02730_),
    .X(_01047_));
 sky130_fd_sc_hd__a31o_1 _20007_ (.A1(_03020_),
    .A2(_03019_),
    .A3(_03025_),
    .B1(\rbzero.pov.spi_done ),
    .X(_03255_));
 sky130_fd_sc_hd__and2_1 _20008_ (.A(_02595_),
    .B(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__clkbuf_1 _20009_ (.A(_03256_),
    .X(_01048_));
 sky130_fd_sc_hd__or4b_1 _20010_ (.A(_04890_),
    .B(_04989_),
    .C(_02703_),
    .D_N(_04990_),
    .X(_03257_));
 sky130_fd_sc_hd__or4bb_1 _20011_ (.A(_04892_),
    .B(_04992_),
    .C_N(_04884_),
    .D_N(_04883_),
    .X(_03258_));
 sky130_fd_sc_hd__inv_2 _20012_ (.A(_04892_),
    .Y(_03259_));
 sky130_fd_sc_hd__or4b_1 _20013_ (.A(_04883_),
    .B(_04992_),
    .C(_03257_),
    .D_N(_04884_),
    .X(_03260_));
 sky130_fd_sc_hd__o21ai_1 _20014_ (.A1(_03259_),
    .A2(_03260_),
    .B1(net71),
    .Y(_03261_));
 sky130_fd_sc_hd__o211a_1 _20015_ (.A1(_03257_),
    .A2(_03258_),
    .B1(_03261_),
    .C1(_03209_),
    .X(_01049_));
 sky130_fd_sc_hd__nor4_1 _20016_ (.A(_03474_),
    .B(_04809_),
    .C(_03554_),
    .D(_04815_),
    .Y(_03262_));
 sky130_fd_sc_hd__or4bb_1 _20017_ (.A(_04006_),
    .B(_04811_),
    .C_N(_04813_),
    .D_N(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__a41o_1 _20018_ (.A1(_04006_),
    .A2(_04811_),
    .A3(_04813_),
    .A4(_03262_),
    .B1(_03911_),
    .X(_03264_));
 sky130_fd_sc_hd__a21oi_1 _20019_ (.A1(net59),
    .A2(_03263_),
    .B1(_03264_),
    .Y(_01050_));
 sky130_fd_sc_hd__or4b_1 _20020_ (.A(_04891_),
    .B(_04887_),
    .C(_04886_),
    .D_N(_04890_),
    .X(_03265_));
 sky130_fd_sc_hd__or4_1 _20021_ (.A(_04990_),
    .B(_04989_),
    .C(_03258_),
    .D(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__and3_1 _20022_ (.A(_04021_),
    .B(_04026_),
    .C(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__nand2_1 _20023_ (.A(_04992_),
    .B(_04037_),
    .Y(_03268_));
 sky130_fd_sc_hd__o211a_1 _20024_ (.A1(_04992_),
    .A2(_03267_),
    .B1(_03268_),
    .C1(_03209_),
    .X(_01051_));
 sky130_fd_sc_hd__a31o_1 _20025_ (.A1(_04892_),
    .A2(_04992_),
    .A3(_04037_),
    .B1(_03911_),
    .X(_03269_));
 sky130_fd_sc_hd__a21oi_1 _20026_ (.A1(_03259_),
    .A2(_03268_),
    .B1(_03269_),
    .Y(_01052_));
 sky130_fd_sc_hd__a21oi_1 _20027_ (.A1(_04892_),
    .A2(_04992_),
    .B1(_04883_),
    .Y(_03270_));
 sky130_fd_sc_hd__nor2_1 _20028_ (.A(_02704_),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__buf_4 _20029_ (.A(_09749_),
    .X(_03272_));
 sky130_fd_sc_hd__a32o_1 _20030_ (.A1(_09753_),
    .A2(_03267_),
    .A3(_03271_),
    .B1(_03272_),
    .B2(_04883_),
    .X(_01053_));
 sky130_fd_sc_hd__nor2_1 _20031_ (.A(_04884_),
    .B(_02704_),
    .Y(_03273_));
 sky130_fd_sc_hd__nor2_1 _20032_ (.A(_02705_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__a32o_1 _20033_ (.A1(_09753_),
    .A2(_03267_),
    .A3(_03274_),
    .B1(_03272_),
    .B2(_04884_),
    .X(_01054_));
 sky130_fd_sc_hd__and3_1 _20034_ (.A(_04989_),
    .B(_04037_),
    .C(_02705_),
    .X(_03275_));
 sky130_fd_sc_hd__a31o_1 _20035_ (.A1(_04021_),
    .A2(_04026_),
    .A3(_02705_),
    .B1(_04989_),
    .X(_03276_));
 sky130_fd_sc_hd__and3b_1 _20036_ (.A_N(_03275_),
    .B(_03276_),
    .C(_05190_),
    .X(_03277_));
 sky130_fd_sc_hd__clkbuf_1 _20037_ (.A(_03277_),
    .X(_01055_));
 sky130_fd_sc_hd__and4_1 _20038_ (.A(_04990_),
    .B(_04989_),
    .C(_04037_),
    .D(_02705_),
    .X(_03278_));
 sky130_fd_sc_hd__nor2_1 _20039_ (.A(_02741_),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__o21a_1 _20040_ (.A1(_04990_),
    .A2(_03275_),
    .B1(_03279_),
    .X(_01056_));
 sky130_fd_sc_hd__a31o_1 _20041_ (.A1(_04886_),
    .A2(_04990_),
    .A3(_03275_),
    .B1(_03911_),
    .X(_03280_));
 sky130_fd_sc_hd__o21ba_1 _20042_ (.A1(_04886_),
    .A2(_03278_),
    .B1_N(_03280_),
    .X(_01057_));
 sky130_fd_sc_hd__and3_1 _20043_ (.A(_04887_),
    .B(_04886_),
    .C(_03278_),
    .X(_03281_));
 sky130_fd_sc_hd__a21o_1 _20044_ (.A1(_04886_),
    .A2(_03278_),
    .B1(_04887_),
    .X(_03282_));
 sky130_fd_sc_hd__and3b_1 _20045_ (.A_N(_03281_),
    .B(_05190_),
    .C(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__clkbuf_1 _20046_ (.A(_03283_),
    .X(_01058_));
 sky130_fd_sc_hd__a31o_1 _20047_ (.A1(_04990_),
    .A2(_04322_),
    .A3(_03275_),
    .B1(_03911_),
    .X(_03284_));
 sky130_fd_sc_hd__o21ba_1 _20048_ (.A1(_04891_),
    .A2(_03281_),
    .B1_N(_03284_),
    .X(_01059_));
 sky130_fd_sc_hd__a21oi_1 _20049_ (.A1(_04891_),
    .A2(_03281_),
    .B1(_04890_),
    .Y(_03285_));
 sky130_fd_sc_hd__inv_2 _20050_ (.A(_03266_),
    .Y(_03286_));
 sky130_fd_sc_hd__a41o_1 _20051_ (.A1(_04990_),
    .A2(_04989_),
    .A3(_04322_),
    .A4(_02705_),
    .B1(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__a31o_1 _20052_ (.A1(_04890_),
    .A2(_04037_),
    .A3(_03287_),
    .B1(_03911_),
    .X(_03288_));
 sky130_fd_sc_hd__nor2_1 _20053_ (.A(_03285_),
    .B(_03288_),
    .Y(_01060_));
 sky130_fd_sc_hd__a31o_1 _20054_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_09753_),
    .A3(_02728_),
    .B1(_02555_),
    .X(_01061_));
 sky130_fd_sc_hd__inv_2 _20056__94 (.A(clknet_1_1__leaf__03045_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _20057__95 (.A(clknet_1_1__leaf__03045_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _20058__96 (.A(clknet_1_1__leaf__03045_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _20059__97 (.A(clknet_1_0__leaf__03045_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _20060__98 (.A(clknet_1_0__leaf__03045_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _20062__99 (.A(clknet_1_1__leaf__03289_),
    .Y(net220));
 sky130_fd_sc_hd__buf_1 _20061_ (.A(clknet_1_0__leaf__03044_),
    .X(_03289_));
 sky130_fd_sc_hd__inv_2 _20063__100 (.A(clknet_1_1__leaf__03289_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _20064__101 (.A(clknet_1_1__leaf__03289_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _20065__102 (.A(clknet_1_1__leaf__03289_),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _20066__103 (.A(clknet_1_1__leaf__03289_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _20067__104 (.A(clknet_1_1__leaf__03289_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _20068__105 (.A(clknet_1_0__leaf__03289_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _20069__106 (.A(clknet_1_0__leaf__03289_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _20070__107 (.A(clknet_1_0__leaf__03289_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _20071__108 (.A(clknet_1_0__leaf__03289_),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _20073__109 (.A(clknet_1_0__leaf__03290_),
    .Y(net230));
 sky130_fd_sc_hd__buf_1 _20072_ (.A(clknet_1_0__leaf__03044_),
    .X(_03290_));
 sky130_fd_sc_hd__inv_2 _20074__110 (.A(clknet_1_0__leaf__03290_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _20075__111 (.A(clknet_1_0__leaf__03290_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _20076__112 (.A(clknet_1_1__leaf__03290_),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _20077__113 (.A(clknet_1_1__leaf__03290_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _20078__114 (.A(clknet_1_1__leaf__03290_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _20079__115 (.A(clknet_1_1__leaf__03290_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20080__116 (.A(clknet_1_1__leaf__03290_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20081__117 (.A(clknet_1_0__leaf__03290_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _20082__118 (.A(clknet_1_0__leaf__03290_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20084__119 (.A(clknet_1_1__leaf__03291_),
    .Y(net240));
 sky130_fd_sc_hd__buf_1 _20083_ (.A(clknet_1_0__leaf__03044_),
    .X(_03291_));
 sky130_fd_sc_hd__inv_2 _20085__120 (.A(clknet_1_1__leaf__03291_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _20086__121 (.A(clknet_1_1__leaf__03291_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20087__122 (.A(clknet_1_1__leaf__03291_),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _20088__123 (.A(clknet_1_1__leaf__03291_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _20089__124 (.A(clknet_1_1__leaf__03291_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _20090__125 (.A(clknet_1_0__leaf__03291_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20091__126 (.A(clknet_1_0__leaf__03291_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20092__127 (.A(clknet_1_0__leaf__03291_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _20093__128 (.A(clknet_1_0__leaf__03291_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20095__129 (.A(clknet_1_0__leaf__03292_),
    .Y(net250));
 sky130_fd_sc_hd__buf_1 _20094_ (.A(clknet_1_0__leaf__03044_),
    .X(_03292_));
 sky130_fd_sc_hd__inv_2 _20096__130 (.A(clknet_1_0__leaf__03292_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _20097__131 (.A(clknet_1_0__leaf__03292_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20098__132 (.A(clknet_1_0__leaf__03292_),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _20099__133 (.A(clknet_1_0__leaf__03292_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _20100__134 (.A(clknet_1_1__leaf__03292_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _20101__135 (.A(clknet_1_1__leaf__03292_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20102__136 (.A(clknet_1_1__leaf__03292_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20103__137 (.A(clknet_1_0__leaf__03292_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _20104__138 (.A(clknet_1_1__leaf__03292_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20106__139 (.A(clknet_1_1__leaf__03293_),
    .Y(net260));
 sky130_fd_sc_hd__buf_1 _20105_ (.A(clknet_1_1__leaf__03044_),
    .X(_03293_));
 sky130_fd_sc_hd__inv_2 _20107__140 (.A(clknet_1_0__leaf__03293_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _20108__141 (.A(clknet_1_0__leaf__03293_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20109__142 (.A(clknet_1_0__leaf__03293_),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _20110__143 (.A(clknet_1_0__leaf__03293_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _20111__144 (.A(clknet_1_0__leaf__03293_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _20112__145 (.A(clknet_1_1__leaf__03293_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20113__146 (.A(clknet_1_1__leaf__03293_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20114__147 (.A(clknet_1_1__leaf__03293_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _20115__148 (.A(clknet_1_1__leaf__03293_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20117__149 (.A(clknet_1_0__leaf__03294_),
    .Y(net270));
 sky130_fd_sc_hd__buf_1 _20116_ (.A(clknet_1_1__leaf__03044_),
    .X(_03294_));
 sky130_fd_sc_hd__inv_2 _20118__150 (.A(clknet_1_0__leaf__03294_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _20119__151 (.A(clknet_1_0__leaf__03294_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20120__152 (.A(clknet_1_0__leaf__03294_),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _20121__153 (.A(clknet_1_0__leaf__03294_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _20122__154 (.A(clknet_1_1__leaf__03294_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _20123__155 (.A(clknet_1_1__leaf__03294_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20124__156 (.A(clknet_1_1__leaf__03294_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20125__157 (.A(clknet_1_1__leaf__03294_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _20126__158 (.A(clknet_1_1__leaf__03294_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20128__159 (.A(clknet_1_1__leaf__03295_),
    .Y(net280));
 sky130_fd_sc_hd__buf_1 _20127_ (.A(clknet_1_0__leaf__03044_),
    .X(_03295_));
 sky130_fd_sc_hd__inv_2 _20129__160 (.A(clknet_1_1__leaf__03295_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _20130__161 (.A(clknet_1_1__leaf__03295_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20131__162 (.A(clknet_1_1__leaf__03295_),
    .Y(net283));
 sky130_fd_sc_hd__inv_2 _20132__163 (.A(clknet_1_1__leaf__03295_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _20133__164 (.A(clknet_1_1__leaf__03295_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _20134__165 (.A(clknet_1_0__leaf__03295_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20135__166 (.A(clknet_1_0__leaf__03295_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20136__167 (.A(clknet_1_0__leaf__03295_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _20137__168 (.A(clknet_1_0__leaf__03295_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20139__169 (.A(clknet_1_0__leaf__03296_),
    .Y(net290));
 sky130_fd_sc_hd__buf_1 _20138_ (.A(clknet_1_0__leaf__03044_),
    .X(_03296_));
 sky130_fd_sc_hd__inv_2 _20140__170 (.A(clknet_1_0__leaf__03296_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _20141__171 (.A(clknet_1_1__leaf__03296_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20142__172 (.A(clknet_1_1__leaf__03296_),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _20143__173 (.A(clknet_1_0__leaf__03296_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _20144__174 (.A(clknet_1_0__leaf__03296_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _20145__175 (.A(clknet_1_0__leaf__03296_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20146__176 (.A(clknet_1_1__leaf__03296_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20147__177 (.A(clknet_1_1__leaf__03296_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _20148__178 (.A(clknet_1_1__leaf__03296_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20150__179 (.A(clknet_1_0__leaf__03297_),
    .Y(net300));
 sky130_fd_sc_hd__buf_1 _20149_ (.A(clknet_1_1__leaf__03044_),
    .X(_03297_));
 sky130_fd_sc_hd__inv_2 _20151__180 (.A(clknet_1_0__leaf__03297_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _20152__181 (.A(clknet_1_0__leaf__03297_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20153__182 (.A(clknet_1_0__leaf__03297_),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _20154__183 (.A(clknet_1_0__leaf__03297_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _20155__184 (.A(clknet_1_0__leaf__03297_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _20156__185 (.A(clknet_1_1__leaf__03297_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20157__186 (.A(clknet_1_1__leaf__03297_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20158__187 (.A(clknet_1_1__leaf__03297_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _20159__188 (.A(clknet_1_1__leaf__03297_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20162__189 (.A(clknet_1_0__leaf__03299_),
    .Y(net310));
 sky130_fd_sc_hd__buf_1 _20160_ (.A(clknet_1_0__leaf__04835_),
    .X(_03298_));
 sky130_fd_sc_hd__buf_1 _20161_ (.A(clknet_1_1__leaf__03298_),
    .X(_03299_));
 sky130_fd_sc_hd__inv_2 _20163__190 (.A(clknet_1_0__leaf__03299_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _20164__191 (.A(clknet_1_0__leaf__03299_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20165__192 (.A(clknet_1_0__leaf__03299_),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 _20166__193 (.A(clknet_1_1__leaf__03299_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _20167__194 (.A(clknet_1_0__leaf__03299_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _20168__195 (.A(clknet_1_0__leaf__03299_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20169__196 (.A(clknet_1_1__leaf__03299_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20170__197 (.A(clknet_1_1__leaf__03299_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _20171__198 (.A(clknet_1_1__leaf__03299_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20173__199 (.A(clknet_1_1__leaf__03300_),
    .Y(net320));
 sky130_fd_sc_hd__buf_1 _20172_ (.A(clknet_1_1__leaf__03298_),
    .X(_03300_));
 sky130_fd_sc_hd__inv_2 _20174__200 (.A(clknet_1_1__leaf__03300_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _20175__201 (.A(clknet_1_1__leaf__03300_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20176__202 (.A(clknet_1_1__leaf__03300_),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _20177__203 (.A(clknet_1_0__leaf__03300_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _20178__204 (.A(clknet_1_1__leaf__03300_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _20179__205 (.A(clknet_1_0__leaf__03300_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20180__206 (.A(clknet_1_0__leaf__03300_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20181__207 (.A(clknet_1_0__leaf__03300_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _20182__208 (.A(clknet_1_0__leaf__03300_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20184__209 (.A(clknet_1_1__leaf__03301_),
    .Y(net330));
 sky130_fd_sc_hd__buf_1 _20183_ (.A(clknet_1_0__leaf__03298_),
    .X(_03301_));
 sky130_fd_sc_hd__inv_2 _20185__210 (.A(clknet_1_1__leaf__03301_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _20186__211 (.A(clknet_1_1__leaf__03301_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20187__212 (.A(clknet_1_0__leaf__03301_),
    .Y(net333));
 sky130_fd_sc_hd__inv_2 _20188__213 (.A(clknet_1_0__leaf__03301_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _20189__214 (.A(clknet_1_0__leaf__03301_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _20190__215 (.A(clknet_1_0__leaf__03301_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20191__216 (.A(clknet_1_1__leaf__03301_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20192__217 (.A(clknet_1_1__leaf__03301_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _20193__218 (.A(clknet_1_1__leaf__03301_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20195__219 (.A(clknet_1_1__leaf__03302_),
    .Y(net340));
 sky130_fd_sc_hd__buf_1 _20194_ (.A(clknet_1_0__leaf__03298_),
    .X(_03302_));
 sky130_fd_sc_hd__inv_2 _20196__220 (.A(clknet_1_1__leaf__03302_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _20197__221 (.A(clknet_1_0__leaf__03302_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20198__222 (.A(clknet_1_0__leaf__03302_),
    .Y(net343));
 sky130_fd_sc_hd__inv_2 _20199__223 (.A(clknet_1_0__leaf__03302_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _20200__224 (.A(clknet_1_0__leaf__03302_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _20201__225 (.A(clknet_1_1__leaf__03302_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20202__226 (.A(clknet_1_1__leaf__03302_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20203__227 (.A(clknet_1_1__leaf__03302_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _20204__228 (.A(clknet_1_1__leaf__03302_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20206__229 (.A(clknet_1_0__leaf__03303_),
    .Y(net350));
 sky130_fd_sc_hd__buf_1 _20205_ (.A(clknet_1_0__leaf__03298_),
    .X(_03303_));
 sky130_fd_sc_hd__inv_2 _20207__230 (.A(clknet_1_0__leaf__03303_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _20208__231 (.A(clknet_1_0__leaf__03303_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20209__232 (.A(clknet_1_0__leaf__03303_),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _20210__233 (.A(clknet_1_1__leaf__03303_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _20211__234 (.A(clknet_1_1__leaf__03303_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _20212__235 (.A(clknet_1_1__leaf__03303_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20213__236 (.A(clknet_1_1__leaf__03303_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20214__237 (.A(clknet_1_1__leaf__03303_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _20215__238 (.A(clknet_1_1__leaf__03303_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20217__239 (.A(clknet_1_0__leaf__03304_),
    .Y(net360));
 sky130_fd_sc_hd__buf_1 _20216_ (.A(clknet_1_1__leaf__03298_),
    .X(_03304_));
 sky130_fd_sc_hd__inv_2 _20218__240 (.A(clknet_1_0__leaf__03304_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _20219__241 (.A(clknet_1_1__leaf__03304_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20220__242 (.A(clknet_1_1__leaf__03304_),
    .Y(net363));
 sky130_fd_sc_hd__inv_2 _20221__243 (.A(clknet_1_1__leaf__03304_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _20222__244 (.A(clknet_1_1__leaf__03304_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _20223__245 (.A(clknet_1_1__leaf__03304_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20224__246 (.A(clknet_1_1__leaf__03304_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20225__247 (.A(clknet_1_0__leaf__03304_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _20226__248 (.A(clknet_1_0__leaf__03304_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20228__249 (.A(clknet_1_0__leaf__03305_),
    .Y(net370));
 sky130_fd_sc_hd__buf_1 _20227_ (.A(clknet_1_1__leaf__03298_),
    .X(_03305_));
 sky130_fd_sc_hd__inv_2 _20229__250 (.A(clknet_1_1__leaf__03305_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _20230__251 (.A(clknet_1_0__leaf__03305_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20231__252 (.A(clknet_1_1__leaf__03305_),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _20232__253 (.A(clknet_1_1__leaf__03305_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _20233__254 (.A(clknet_1_0__leaf__03305_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _20234__255 (.A(clknet_1_0__leaf__03305_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20235__256 (.A(clknet_1_1__leaf__03305_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20236__257 (.A(clknet_1_1__leaf__03305_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _20237__258 (.A(clknet_1_1__leaf__03305_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20239__259 (.A(clknet_1_0__leaf__03306_),
    .Y(net380));
 sky130_fd_sc_hd__buf_1 _20238_ (.A(clknet_1_0__leaf__03298_),
    .X(_03306_));
 sky130_fd_sc_hd__inv_2 _20240__260 (.A(clknet_1_1__leaf__03306_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _20241__261 (.A(clknet_1_1__leaf__03306_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20242__262 (.A(clknet_1_1__leaf__03306_),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _20243__263 (.A(clknet_1_1__leaf__03306_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _20244__264 (.A(clknet_1_0__leaf__03306_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _20245__265 (.A(clknet_1_1__leaf__03306_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20246__266 (.A(clknet_1_1__leaf__03306_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20247__267 (.A(clknet_1_0__leaf__03306_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _20248__268 (.A(clknet_1_0__leaf__03306_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20250__269 (.A(clknet_1_1__leaf__03307_),
    .Y(net390));
 sky130_fd_sc_hd__buf_1 _20249_ (.A(clknet_1_0__leaf__03298_),
    .X(_03307_));
 sky130_fd_sc_hd__inv_2 _20251__270 (.A(clknet_1_1__leaf__03307_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _20252__271 (.A(clknet_1_1__leaf__03307_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20253__272 (.A(clknet_1_1__leaf__03307_),
    .Y(net393));
 sky130_fd_sc_hd__inv_2 _20254__273 (.A(clknet_1_0__leaf__03307_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _20255__274 (.A(clknet_1_1__leaf__03307_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _20256__275 (.A(clknet_1_0__leaf__03307_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20257__276 (.A(clknet_1_0__leaf__03307_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20258__277 (.A(clknet_1_0__leaf__03307_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _20259__278 (.A(clknet_1_0__leaf__03307_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20261__279 (.A(clknet_1_0__leaf__03308_),
    .Y(net400));
 sky130_fd_sc_hd__buf_1 _20260_ (.A(clknet_1_0__leaf__03298_),
    .X(_03308_));
 sky130_fd_sc_hd__inv_2 _20262__280 (.A(clknet_1_0__leaf__03308_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _20263__281 (.A(clknet_1_0__leaf__03308_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20264__282 (.A(clknet_1_0__leaf__03308_),
    .Y(net403));
 sky130_fd_sc_hd__inv_2 _20265__283 (.A(clknet_1_1__leaf__03308_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _20266__284 (.A(clknet_1_0__leaf__03308_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _20267__285 (.A(clknet_1_1__leaf__03308_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20268__286 (.A(clknet_1_1__leaf__03308_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20269__287 (.A(clknet_1_1__leaf__03308_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _20270__288 (.A(clknet_1_1__leaf__03308_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20273__289 (.A(clknet_1_1__leaf__03310_),
    .Y(net410));
 sky130_fd_sc_hd__buf_1 _20271_ (.A(clknet_1_0__leaf__04835_),
    .X(_03309_));
 sky130_fd_sc_hd__buf_1 _20272_ (.A(clknet_1_1__leaf__03309_),
    .X(_03310_));
 sky130_fd_sc_hd__inv_2 _20274__290 (.A(clknet_1_1__leaf__03310_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _20275__291 (.A(clknet_1_1__leaf__03310_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20276__292 (.A(clknet_1_1__leaf__03310_),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _20277__293 (.A(clknet_1_0__leaf__03310_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _20278__294 (.A(clknet_1_0__leaf__03310_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _20279__295 (.A(clknet_1_0__leaf__03310_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20280__296 (.A(clknet_1_1__leaf__03310_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20281__297 (.A(clknet_1_0__leaf__03310_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _20282__298 (.A(clknet_1_0__leaf__03310_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20284__299 (.A(clknet_1_0__leaf__03311_),
    .Y(net420));
 sky130_fd_sc_hd__buf_1 _20283_ (.A(clknet_1_1__leaf__03309_),
    .X(_03311_));
 sky130_fd_sc_hd__inv_2 _20285__300 (.A(clknet_1_0__leaf__03311_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _20286__301 (.A(clknet_1_0__leaf__03311_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20287__302 (.A(clknet_1_0__leaf__03311_),
    .Y(net423));
 sky130_fd_sc_hd__inv_2 _20288__303 (.A(clknet_1_0__leaf__03311_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _20289__304 (.A(clknet_1_0__leaf__03311_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _20290__305 (.A(clknet_1_1__leaf__03311_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20291__306 (.A(clknet_1_1__leaf__03311_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20292__307 (.A(clknet_1_1__leaf__03311_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _20293__308 (.A(clknet_1_1__leaf__03311_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20295__309 (.A(clknet_1_0__leaf__03312_),
    .Y(net430));
 sky130_fd_sc_hd__buf_1 _20294_ (.A(clknet_1_1__leaf__03309_),
    .X(_03312_));
 sky130_fd_sc_hd__inv_2 _20296__310 (.A(clknet_1_0__leaf__03312_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _20297__311 (.A(clknet_1_0__leaf__03312_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20298__312 (.A(clknet_1_1__leaf__03312_),
    .Y(net433));
 sky130_fd_sc_hd__inv_2 _20299__313 (.A(clknet_1_1__leaf__03312_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _20300__314 (.A(clknet_1_1__leaf__03312_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _20301__315 (.A(clknet_1_1__leaf__03312_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20302__316 (.A(clknet_1_0__leaf__03312_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20303__317 (.A(clknet_1_0__leaf__03312_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _20304__318 (.A(clknet_1_0__leaf__03312_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20306__319 (.A(clknet_1_1__leaf__03313_),
    .Y(net440));
 sky130_fd_sc_hd__buf_1 _20305_ (.A(clknet_1_1__leaf__03309_),
    .X(_03313_));
 sky130_fd_sc_hd__inv_2 _20307__320 (.A(clknet_1_1__leaf__03313_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _20308__321 (.A(clknet_1_0__leaf__03313_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20309__322 (.A(clknet_1_0__leaf__03313_),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 _20310__323 (.A(clknet_1_0__leaf__03313_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _20311__324 (.A(clknet_1_0__leaf__03313_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _20312__325 (.A(clknet_1_1__leaf__03313_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20313__326 (.A(clknet_1_1__leaf__03313_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20314__327 (.A(clknet_1_1__leaf__03313_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _20315__328 (.A(clknet_1_0__leaf__03313_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20317__329 (.A(clknet_1_0__leaf__03314_),
    .Y(net450));
 sky130_fd_sc_hd__buf_1 _20316_ (.A(clknet_1_1__leaf__03309_),
    .X(_03314_));
 sky130_fd_sc_hd__inv_2 _20318__330 (.A(clknet_1_0__leaf__03314_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _20319__331 (.A(clknet_1_0__leaf__03314_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20320__332 (.A(clknet_1_0__leaf__03314_),
    .Y(net453));
 sky130_fd_sc_hd__inv_2 _20321__333 (.A(clknet_1_1__leaf__03314_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _20322__334 (.A(clknet_1_1__leaf__03314_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _20323__335 (.A(clknet_1_1__leaf__03314_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20324__336 (.A(clknet_1_1__leaf__03314_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20325__337 (.A(clknet_1_1__leaf__03314_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _20326__338 (.A(clknet_1_1__leaf__03314_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20328__339 (.A(clknet_1_0__leaf__03315_),
    .Y(net460));
 sky130_fd_sc_hd__buf_1 _20327_ (.A(clknet_1_1__leaf__03309_),
    .X(_03315_));
 sky130_fd_sc_hd__inv_2 _20329__340 (.A(clknet_1_0__leaf__03315_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _20330__341 (.A(clknet_1_0__leaf__03315_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20331__342 (.A(clknet_1_0__leaf__03315_),
    .Y(net463));
 sky130_fd_sc_hd__inv_2 _20332__343 (.A(clknet_1_1__leaf__03315_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _20333__344 (.A(clknet_1_1__leaf__03315_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _20334__345 (.A(clknet_1_1__leaf__03315_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20335__346 (.A(clknet_1_1__leaf__03315_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20336__347 (.A(clknet_1_1__leaf__03315_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _20337__348 (.A(clknet_1_0__leaf__03315_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20339__349 (.A(clknet_1_1__leaf__03316_),
    .Y(net470));
 sky130_fd_sc_hd__buf_1 _20338_ (.A(clknet_1_0__leaf__03309_),
    .X(_03316_));
 sky130_fd_sc_hd__inv_2 _20340__350 (.A(clknet_1_1__leaf__03316_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _20341__351 (.A(clknet_1_1__leaf__03316_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20342__352 (.A(clknet_1_1__leaf__03316_),
    .Y(net473));
 sky130_fd_sc_hd__inv_2 _20343__353 (.A(clknet_1_0__leaf__03316_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _20344__354 (.A(clknet_1_0__leaf__03316_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _20345__355 (.A(clknet_1_0__leaf__03316_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20346__356 (.A(clknet_1_0__leaf__03316_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20347__357 (.A(clknet_1_0__leaf__03316_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _20348__358 (.A(clknet_1_1__leaf__03316_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20350__359 (.A(clknet_1_0__leaf__03317_),
    .Y(net480));
 sky130_fd_sc_hd__buf_1 _20349_ (.A(clknet_1_0__leaf__03309_),
    .X(_03317_));
 sky130_fd_sc_hd__inv_2 _20351__360 (.A(clknet_1_0__leaf__03317_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _20352__361 (.A(clknet_1_0__leaf__03317_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20353__362 (.A(clknet_1_0__leaf__03317_),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _20354__363 (.A(clknet_1_0__leaf__03317_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _20355__364 (.A(clknet_1_0__leaf__03317_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _20356__365 (.A(clknet_1_1__leaf__03317_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20357__366 (.A(clknet_1_1__leaf__03317_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20358__367 (.A(clknet_1_1__leaf__03317_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _20359__368 (.A(clknet_1_1__leaf__03317_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20361__369 (.A(clknet_1_0__leaf__03318_),
    .Y(net490));
 sky130_fd_sc_hd__buf_1 _20360_ (.A(clknet_1_0__leaf__03309_),
    .X(_03318_));
 sky130_fd_sc_hd__inv_2 _20362__370 (.A(clknet_1_0__leaf__03318_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _20363__371 (.A(clknet_1_0__leaf__03318_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20364__372 (.A(clknet_1_0__leaf__03318_),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _20365__373 (.A(clknet_1_1__leaf__03318_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _20366__374 (.A(clknet_1_1__leaf__03318_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _20367__375 (.A(clknet_1_1__leaf__03318_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20368__376 (.A(clknet_1_1__leaf__03318_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20369__377 (.A(clknet_1_1__leaf__03318_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _20370__378 (.A(clknet_1_0__leaf__03318_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20372__379 (.A(clknet_1_0__leaf__03319_),
    .Y(net500));
 sky130_fd_sc_hd__buf_1 _20371_ (.A(clknet_1_0__leaf__03309_),
    .X(_03319_));
 sky130_fd_sc_hd__inv_2 _20373__380 (.A(clknet_1_0__leaf__03319_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _20374__381 (.A(clknet_1_0__leaf__03319_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20375__382 (.A(clknet_1_0__leaf__03319_),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _20376__383 (.A(clknet_1_0__leaf__03319_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _20377__384 (.A(clknet_1_0__leaf__03319_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _20378__385 (.A(clknet_1_1__leaf__03319_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20379__386 (.A(clknet_1_1__leaf__03319_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20380__387 (.A(clknet_1_1__leaf__03319_),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _20381__388 (.A(clknet_1_1__leaf__03319_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _12189__389 (.A(_04959_),
    .Y(net510));
 sky130_fd_sc_hd__buf_1 _20382_ (.A(clknet_1_0__leaf__04835_),
    .X(_03320_));
 sky130_fd_sc_hd__inv_2 _20384__10 (.A(clknet_1_0__leaf__03320_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _20385__11 (.A(clknet_1_0__leaf__03320_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _20386__12 (.A(clknet_1_0__leaf__03320_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _20387__13 (.A(clknet_1_1__leaf__03320_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _20388__14 (.A(clknet_1_1__leaf__03320_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _20389__15 (.A(clknet_1_1__leaf__03320_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _20390__16 (.A(clknet_1_1__leaf__03320_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _20391__17 (.A(clknet_1_0__leaf__03320_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _20392__18 (.A(clknet_1_0__leaf__03320_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _20394__19 (.A(clknet_1_1__leaf__03321_),
    .Y(net140));
 sky130_fd_sc_hd__buf_1 _20393_ (.A(clknet_1_0__leaf__04835_),
    .X(_03321_));
 sky130_fd_sc_hd__inv_2 _20395__20 (.A(clknet_1_1__leaf__03321_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _20396__21 (.A(clknet_1_1__leaf__03321_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _20397__22 (.A(clknet_1_1__leaf__03321_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _20398__23 (.A(clknet_1_0__leaf__03321_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _20399__24 (.A(clknet_1_0__leaf__03321_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _20400__25 (.A(clknet_1_0__leaf__03321_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20401__26 (.A(clknet_1_0__leaf__03321_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20402__27 (.A(clknet_1_1__leaf__03321_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _20403__28 (.A(clknet_1_0__leaf__03321_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _19572__29 (.A(clknet_1_1__leaf__03038_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _20405__6 (.A(clknet_1_1__leaf__03037_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _20406__7 (.A(clknet_1_1__leaf__03037_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _20407__8 (.A(clknet_1_1__leaf__03037_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _20383__9 (.A(clknet_1_0__leaf__03320_),
    .Y(net130));
 sky130_fd_sc_hd__nor2_1 _20408_ (.A(\gpout5.clk_div[0] ),
    .B(net60),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2_1 _20409_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_03322_));
 sky130_fd_sc_hd__or2_1 _20410_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_03323_));
 sky130_fd_sc_hd__and3_1 _20411_ (.A(_02721_),
    .B(_03322_),
    .C(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_1 _20412_ (.A(_03324_),
    .X(_01383_));
 sky130_fd_sc_hd__nand2_1 _20413_ (.A(\rbzero.traced_texa[-12] ),
    .B(\rbzero.texV[-12] ),
    .Y(_03325_));
 sky130_fd_sc_hd__or2_1 _20414_ (.A(\rbzero.traced_texa[-12] ),
    .B(\rbzero.texV[-12] ),
    .X(_03326_));
 sky130_fd_sc_hd__buf_4 _20415_ (.A(_02695_),
    .X(_03327_));
 sky130_fd_sc_hd__a32o_1 _20416_ (.A1(_03272_),
    .A2(_03325_),
    .A3(_03326_),
    .B1(_03327_),
    .B2(\rbzero.texV[-12] ),
    .X(_01384_));
 sky130_fd_sc_hd__or2_1 _20417_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_03328_));
 sky130_fd_sc_hd__nand2_1 _20418_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_03329_));
 sky130_fd_sc_hd__nand3b_1 _20419_ (.A_N(_03325_),
    .B(_03328_),
    .C(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__a21bo_1 _20420_ (.A1(_03328_),
    .A2(_03329_),
    .B1_N(_03325_),
    .X(_03331_));
 sky130_fd_sc_hd__a32o_1 _20421_ (.A1(_03272_),
    .A2(_03330_),
    .A3(_03331_),
    .B1(_03327_),
    .B2(\rbzero.texV[-11] ),
    .X(_01385_));
 sky130_fd_sc_hd__clkbuf_4 _20422_ (.A(_09750_),
    .X(_03332_));
 sky130_fd_sc_hd__and2_1 _20423_ (.A(_03329_),
    .B(_03330_),
    .X(_03333_));
 sky130_fd_sc_hd__nor2_1 _20424_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03334_));
 sky130_fd_sc_hd__nand2_1 _20425_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03335_));
 sky130_fd_sc_hd__and2b_1 _20426_ (.A_N(_03334_),
    .B(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__xnor2_1 _20427_ (.A(_03333_),
    .B(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__a22o_1 _20428_ (.A1(\rbzero.texV[-10] ),
    .A2(_03175_),
    .B1(_03332_),
    .B2(_03337_),
    .X(_01386_));
 sky130_fd_sc_hd__or2_1 _20429_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .X(_03338_));
 sky130_fd_sc_hd__nand2_1 _20430_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03339_));
 sky130_fd_sc_hd__nand2_1 _20431_ (.A(_03338_),
    .B(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__o21ai_1 _20432_ (.A1(_03333_),
    .A2(_03334_),
    .B1(_03335_),
    .Y(_03341_));
 sky130_fd_sc_hd__xnor2_1 _20433_ (.A(_03340_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__a22o_1 _20434_ (.A1(\rbzero.texV[-9] ),
    .A2(_03175_),
    .B1(_03332_),
    .B2(_03342_),
    .X(_01387_));
 sky130_fd_sc_hd__nor2_1 _20435_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03343_));
 sky130_fd_sc_hd__and2_1 _20436_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .X(_03344_));
 sky130_fd_sc_hd__a21boi_1 _20437_ (.A1(_03338_),
    .A2(_03341_),
    .B1_N(_03339_),
    .Y(_03345_));
 sky130_fd_sc_hd__o21ai_1 _20438_ (.A1(_03343_),
    .A2(_03344_),
    .B1(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__or3_1 _20439_ (.A(_03343_),
    .B(_03344_),
    .C(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__a32o_1 _20440_ (.A1(_03272_),
    .A2(_03346_),
    .A3(_03347_),
    .B1(_03327_),
    .B2(\rbzero.texV[-8] ),
    .X(_01388_));
 sky130_fd_sc_hd__xnor2_1 _20441_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_03348_));
 sky130_fd_sc_hd__o21bai_1 _20442_ (.A1(_03343_),
    .A2(_03345_),
    .B1_N(_03344_),
    .Y(_03349_));
 sky130_fd_sc_hd__xnor2_1 _20443_ (.A(_03348_),
    .B(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__a22o_1 _20444_ (.A1(\rbzero.texV[-7] ),
    .A2(_03175_),
    .B1(_03332_),
    .B2(_03350_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2_1 _20445_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _20446_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03352_));
 sky130_fd_sc_hd__and2b_1 _20447_ (.A_N(_03351_),
    .B(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__a21o_1 _20448_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(\rbzero.texV[-7] ),
    .B1(_03349_),
    .X(_03354_));
 sky130_fd_sc_hd__o21ai_1 _20449_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(\rbzero.texV[-7] ),
    .B1(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__xnor2_1 _20450_ (.A(_03353_),
    .B(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__a22o_1 _20451_ (.A1(\rbzero.texV[-6] ),
    .A2(_03175_),
    .B1(_03332_),
    .B2(_03356_),
    .X(_01390_));
 sky130_fd_sc_hd__or2_1 _20452_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .X(_03357_));
 sky130_fd_sc_hd__nand2_1 _20453_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03358_));
 sky130_fd_sc_hd__o21ai_1 _20454_ (.A1(_03351_),
    .A2(_03355_),
    .B1(_03352_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand3_1 _20455_ (.A(_03357_),
    .B(_03358_),
    .C(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__a21o_1 _20456_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03359_),
    .X(_03361_));
 sky130_fd_sc_hd__a32o_1 _20457_ (.A1(_03272_),
    .A2(_03360_),
    .A3(_03361_),
    .B1(_03327_),
    .B2(\rbzero.texV[-5] ),
    .X(_01391_));
 sky130_fd_sc_hd__nor2_1 _20458_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03362_));
 sky130_fd_sc_hd__and2_1 _20459_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .X(_03363_));
 sky130_fd_sc_hd__a21boi_1 _20460_ (.A1(_03357_),
    .A2(_03359_),
    .B1_N(_03358_),
    .Y(_03364_));
 sky130_fd_sc_hd__or3_1 _20461_ (.A(_03362_),
    .B(_03363_),
    .C(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__o21ai_1 _20462_ (.A1(_03362_),
    .A2(_03363_),
    .B1(_03364_),
    .Y(_03366_));
 sky130_fd_sc_hd__a32o_1 _20463_ (.A1(_03272_),
    .A2(_03365_),
    .A3(_03366_),
    .B1(_03327_),
    .B2(\rbzero.texV[-4] ),
    .X(_01392_));
 sky130_fd_sc_hd__or2_1 _20464_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .X(_03367_));
 sky130_fd_sc_hd__nand2_1 _20465_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03368_));
 sky130_fd_sc_hd__o21bai_1 _20466_ (.A1(_03362_),
    .A2(_03364_),
    .B1_N(_03363_),
    .Y(_03369_));
 sky130_fd_sc_hd__a21o_1 _20467_ (.A1(_03367_),
    .A2(_03368_),
    .B1(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__nand3_1 _20468_ (.A(_03367_),
    .B(_03368_),
    .C(_03369_),
    .Y(_03371_));
 sky130_fd_sc_hd__a32o_1 _20469_ (.A1(_03272_),
    .A2(_03370_),
    .A3(_03371_),
    .B1(_03250_),
    .B2(\rbzero.texV[-3] ),
    .X(_01393_));
 sky130_fd_sc_hd__nor2_1 _20470_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_03372_));
 sky130_fd_sc_hd__and2_1 _20471_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_03373_));
 sky130_fd_sc_hd__or2_1 _20472_ (.A(_03372_),
    .B(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__a21boi_1 _20473_ (.A1(_03367_),
    .A2(_03369_),
    .B1_N(_03368_),
    .Y(_03375_));
 sky130_fd_sc_hd__xor2_1 _20474_ (.A(_03374_),
    .B(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__a22o_1 _20475_ (.A1(\rbzero.texV[-2] ),
    .A2(_03175_),
    .B1(_03332_),
    .B2(_03376_),
    .X(_01394_));
 sky130_fd_sc_hd__nor2_1 _20476_ (.A(_03374_),
    .B(_03375_),
    .Y(_03377_));
 sky130_fd_sc_hd__or2_1 _20477_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_03378_));
 sky130_fd_sc_hd__nand2_1 _20478_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_03379_));
 sky130_fd_sc_hd__o211a_1 _20479_ (.A1(_03373_),
    .A2(_03377_),
    .B1(_03378_),
    .C1(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__inv_2 _20480_ (.A(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__a211o_1 _20481_ (.A1(_03378_),
    .A2(_03379_),
    .B1(_03373_),
    .C1(_03377_),
    .X(_03382_));
 sky130_fd_sc_hd__a32o_1 _20482_ (.A1(_03272_),
    .A2(_03381_),
    .A3(_03382_),
    .B1(_03250_),
    .B2(\rbzero.texV[-1] ),
    .X(_01395_));
 sky130_fd_sc_hd__or2_1 _20483_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_03383_));
 sky130_fd_sc_hd__nand2_1 _20484_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_1 _20485_ (.A(_03379_),
    .B(_03381_),
    .Y(_03385_));
 sky130_fd_sc_hd__a21o_1 _20486_ (.A1(_03383_),
    .A2(_03384_),
    .B1(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__and3_1 _20487_ (.A(_03383_),
    .B(_03384_),
    .C(_03385_),
    .X(_03387_));
 sky130_fd_sc_hd__inv_2 _20488_ (.A(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__a32o_1 _20489_ (.A1(_03272_),
    .A2(_03386_),
    .A3(_03388_),
    .B1(_03250_),
    .B2(\rbzero.texV[0] ),
    .X(_01396_));
 sky130_fd_sc_hd__or2_1 _20490_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_03389_));
 sky130_fd_sc_hd__nand2_1 _20491_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_03390_));
 sky130_fd_sc_hd__nand2_1 _20492_ (.A(_03384_),
    .B(_03388_),
    .Y(_03391_));
 sky130_fd_sc_hd__a21o_1 _20493_ (.A1(_03389_),
    .A2(_03390_),
    .B1(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__and3_1 _20494_ (.A(_03389_),
    .B(_03390_),
    .C(_03391_),
    .X(_03393_));
 sky130_fd_sc_hd__inv_2 _20495_ (.A(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__a32o_1 _20496_ (.A1(_09750_),
    .A2(_03392_),
    .A3(_03394_),
    .B1(_03250_),
    .B2(\rbzero.texV[1] ),
    .X(_01397_));
 sky130_fd_sc_hd__or2_1 _20497_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_03395_));
 sky130_fd_sc_hd__nand2_1 _20498_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_03396_));
 sky130_fd_sc_hd__nand2_1 _20499_ (.A(_03390_),
    .B(_03394_),
    .Y(_03397_));
 sky130_fd_sc_hd__and3_1 _20500_ (.A(_03395_),
    .B(_03396_),
    .C(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__inv_2 _20501_ (.A(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__a21o_1 _20502_ (.A1(_03395_),
    .A2(_03396_),
    .B1(_03397_),
    .X(_03400_));
 sky130_fd_sc_hd__a32o_1 _20503_ (.A1(_09750_),
    .A2(_03399_),
    .A3(_03400_),
    .B1(_03250_),
    .B2(\rbzero.texV[2] ),
    .X(_01398_));
 sky130_fd_sc_hd__or2_1 _20504_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_03401_));
 sky130_fd_sc_hd__nand2_1 _20505_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _20506_ (.A(_03396_),
    .B(_03399_),
    .Y(_03403_));
 sky130_fd_sc_hd__a21o_1 _20507_ (.A1(_03401_),
    .A2(_03402_),
    .B1(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__nand3_1 _20508_ (.A(_03401_),
    .B(_03402_),
    .C(_03403_),
    .Y(_03405_));
 sky130_fd_sc_hd__a32o_1 _20509_ (.A1(_09750_),
    .A2(_03404_),
    .A3(_03405_),
    .B1(_03250_),
    .B2(\rbzero.texV[3] ),
    .X(_01399_));
 sky130_fd_sc_hd__a21boi_1 _20510_ (.A1(_03401_),
    .A2(_03403_),
    .B1_N(_03402_),
    .Y(_03406_));
 sky130_fd_sc_hd__nor2_1 _20511_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _20512_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03408_));
 sky130_fd_sc_hd__and2b_1 _20513_ (.A_N(_03407_),
    .B(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__xnor2_1 _20514_ (.A(_03406_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__a22o_1 _20515_ (.A1(\rbzero.texV[4] ),
    .A2(_03327_),
    .B1(_03332_),
    .B2(_03410_),
    .X(_01400_));
 sky130_fd_sc_hd__or2_1 _20516_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .X(_03411_));
 sky130_fd_sc_hd__nand2_1 _20517_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03412_));
 sky130_fd_sc_hd__nand2_1 _20518_ (.A(_03411_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__o21ai_1 _20519_ (.A1(_03406_),
    .A2(_03407_),
    .B1(_03408_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_1 _20520_ (.A(_03413_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__a22o_1 _20521_ (.A1(\rbzero.texV[5] ),
    .A2(_03327_),
    .B1(_03332_),
    .B2(_03415_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2_1 _20522_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_1 _20523_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03417_));
 sky130_fd_sc_hd__and2b_1 _20524_ (.A_N(_03416_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__a21boi_1 _20525_ (.A1(_03411_),
    .A2(_03414_),
    .B1_N(_03412_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_1 _20526_ (.A(_03418_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__a22o_1 _20527_ (.A1(\rbzero.texV[6] ),
    .A2(_03327_),
    .B1(_03332_),
    .B2(_03420_),
    .X(_01402_));
 sky130_fd_sc_hd__xnor2_1 _20528_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03421_));
 sky130_fd_sc_hd__o21ai_1 _20529_ (.A1(_03416_),
    .A2(_03419_),
    .B1(_03417_),
    .Y(_03422_));
 sky130_fd_sc_hd__xnor2_1 _20530_ (.A(_03421_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__a22o_1 _20531_ (.A1(\rbzero.texV[7] ),
    .A2(_03327_),
    .B1(_03332_),
    .B2(_03423_),
    .X(_01403_));
 sky130_fd_sc_hd__nor2_1 _20532_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03424_));
 sky130_fd_sc_hd__nand2_1 _20533_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03425_));
 sky130_fd_sc_hd__and2b_1 _20534_ (.A_N(_03424_),
    .B(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__a21o_1 _20535_ (.A1(\rbzero.traced_texa[7] ),
    .A2(\rbzero.texV[7] ),
    .B1(_03422_),
    .X(_03427_));
 sky130_fd_sc_hd__o21ai_1 _20536_ (.A1(\rbzero.traced_texa[7] ),
    .A2(\rbzero.texV[7] ),
    .B1(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__xnor2_1 _20537_ (.A(_03426_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__a22o_1 _20538_ (.A1(\rbzero.texV[8] ),
    .A2(_03327_),
    .B1(_03332_),
    .B2(_03429_),
    .X(_01404_));
 sky130_fd_sc_hd__or2_1 _20539_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_1 _20540_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03431_));
 sky130_fd_sc_hd__o21ai_1 _20541_ (.A1(_03424_),
    .A2(_03428_),
    .B1(_03425_),
    .Y(_03432_));
 sky130_fd_sc_hd__a21o_1 _20542_ (.A1(_03430_),
    .A2(_03431_),
    .B1(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__nand3_1 _20543_ (.A(_03430_),
    .B(_03431_),
    .C(_03432_),
    .Y(_03434_));
 sky130_fd_sc_hd__a32o_1 _20544_ (.A1(_09750_),
    .A2(_03433_),
    .A3(_03434_),
    .B1(_03250_),
    .B2(\rbzero.texV[9] ),
    .X(_01405_));
 sky130_fd_sc_hd__or2_1 _20545_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .X(_03435_));
 sky130_fd_sc_hd__nand2_1 _20546_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_03436_));
 sky130_fd_sc_hd__a21o_1 _20547_ (.A1(\rbzero.traced_texa[9] ),
    .A2(\rbzero.texV[9] ),
    .B1(_03432_),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_1 _20548_ (.A1(_03435_),
    .A2(_03436_),
    .B1(_03437_),
    .B2(_03430_),
    .X(_03438_));
 sky130_fd_sc_hd__nand4_1 _20549_ (.A(_03430_),
    .B(_03435_),
    .C(_03436_),
    .D(_03437_),
    .Y(_03439_));
 sky130_fd_sc_hd__a32o_1 _20550_ (.A1(_09750_),
    .A2(_03438_),
    .A3(_03439_),
    .B1(_03250_),
    .B2(\rbzero.texV[10] ),
    .X(_01406_));
 sky130_fd_sc_hd__xnor2_1 _20551_ (.A(\rbzero.traced_texa[11] ),
    .B(\rbzero.texV[11] ),
    .Y(_03440_));
 sky130_fd_sc_hd__a21oi_1 _20552_ (.A1(_03436_),
    .A2(_03439_),
    .B1(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__a31o_1 _20553_ (.A1(_03436_),
    .A2(_03439_),
    .A3(_03440_),
    .B1(_09748_),
    .X(_03442_));
 sky130_fd_sc_hd__a2bb2o_1 _20554_ (.A1_N(_03441_),
    .A2_N(_03442_),
    .B1(\rbzero.texV[11] ),
    .B2(net60),
    .X(_01407_));
 sky130_fd_sc_hd__a22o_1 _20555_ (.A1(\rbzero.traced_texVinit[0] ),
    .A2(_09770_),
    .B1(_09771_),
    .B2(_09068_),
    .X(_01408_));
 sky130_fd_sc_hd__buf_4 _20556_ (.A(_07695_),
    .X(_03443_));
 sky130_fd_sc_hd__a22o_1 _20557_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_03443_),
    .B1(_09771_),
    .B2(_09076_),
    .X(_01409_));
 sky130_fd_sc_hd__a2bb2o_1 _20558_ (.A1_N(_09763_),
    .A2_N(_09859_),
    .B1(\rbzero.traced_texVinit[2] ),
    .B2(_09762_),
    .X(_01410_));
 sky130_fd_sc_hd__a2bb2o_1 _20559_ (.A1_N(_09763_),
    .A2_N(_09194_),
    .B1(\rbzero.traced_texVinit[3] ),
    .B2(_09762_),
    .X(_01411_));
 sky130_fd_sc_hd__inv_2 _20560_ (.A(_09331_),
    .Y(_03444_));
 sky130_fd_sc_hd__a22o_1 _20561_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_03443_),
    .B1(_09771_),
    .B2(_03444_),
    .X(_01412_));
 sky130_fd_sc_hd__a2bb2o_1 _20562_ (.A1_N(_07831_),
    .A2_N(_09458_),
    .B1(\rbzero.traced_texVinit[5] ),
    .B2(_09762_),
    .X(_01413_));
 sky130_fd_sc_hd__a22o_1 _20563_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_03443_),
    .B1(_09771_),
    .B2(_09597_),
    .X(_01414_));
 sky130_fd_sc_hd__a22o_1 _20564_ (.A1(\rbzero.traced_texVinit[7] ),
    .A2(_03443_),
    .B1(_09771_),
    .B2(_09739_),
    .X(_01415_));
 sky130_fd_sc_hd__o2bb2ai_1 _20565_ (.A1_N(\rbzero.traced_texVinit[8] ),
    .A2_N(_09764_),
    .B1(_07831_),
    .B2(_10027_),
    .Y(_01416_));
 sky130_fd_sc_hd__o2bb2ai_1 _20566_ (.A1_N(\rbzero.traced_texVinit[9] ),
    .A2_N(_09764_),
    .B1(_07831_),
    .B2(_10171_),
    .Y(_01417_));
 sky130_fd_sc_hd__a22o_1 _20567_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_03443_),
    .B1(_09771_),
    .B2(_10297_),
    .X(_01418_));
 sky130_fd_sc_hd__a22o_1 _20568_ (.A1(\rbzero.traced_texVinit[11] ),
    .A2(_03443_),
    .B1(_07756_),
    .B2(_01552_),
    .X(_01419_));
 sky130_fd_sc_hd__nor2_1 _20569_ (.A(\gpout0.clk_div[0] ),
    .B(net60),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _20570_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_03445_));
 sky130_fd_sc_hd__or2_1 _20571_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_03446_));
 sky130_fd_sc_hd__and3_1 _20572_ (.A(_02721_),
    .B(_03445_),
    .C(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _20573_ (.A(_03447_),
    .X(_01421_));
 sky130_fd_sc_hd__nor2_1 _20574_ (.A(\gpout1.clk_div[0] ),
    .B(net60),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _20575_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_03448_));
 sky130_fd_sc_hd__or2_1 _20576_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_03449_));
 sky130_fd_sc_hd__and3_1 _20577_ (.A(_02721_),
    .B(_03448_),
    .C(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _20578_ (.A(_03450_),
    .X(_01423_));
 sky130_fd_sc_hd__or2_1 _20579_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_03451_));
 sky130_fd_sc_hd__a32o_1 _20580_ (.A1(_07685_),
    .A2(_07679_),
    .A3(_03451_),
    .B1(_03443_),
    .B2(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_01424_));
 sky130_fd_sc_hd__a21bo_1 _20581_ (.A1(_07687_),
    .A2(_07686_),
    .B1_N(_07685_),
    .X(_03452_));
 sky130_fd_sc_hd__nor2_1 _20582_ (.A(_07688_),
    .B(_07831_),
    .Y(_03453_));
 sky130_fd_sc_hd__a22o_1 _20583_ (.A1(\rbzero.wall_tracer.rayAddendX[-8] ),
    .A2(_03443_),
    .B1(_03452_),
    .B2(_03453_),
    .X(_01425_));
 sky130_fd_sc_hd__and2b_1 _20584_ (.A_N(_07684_),
    .B(_07690_),
    .X(_03454_));
 sky130_fd_sc_hd__xnor2_1 _20585_ (.A(_07689_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__a22o_1 _20586_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_03443_),
    .B1(_07756_),
    .B2(_03455_),
    .X(_01426_));
 sky130_fd_sc_hd__a21oi_1 _20587_ (.A1(_07683_),
    .A2(_07692_),
    .B1(_07691_),
    .Y(_03456_));
 sky130_fd_sc_hd__a31o_1 _20588_ (.A1(_07683_),
    .A2(_07692_),
    .A3(_07691_),
    .B1(_07831_),
    .X(_03457_));
 sky130_fd_sc_hd__a2bb2o_1 _20589_ (.A1_N(_03456_),
    .A2_N(_03457_),
    .B1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B2(_09762_),
    .X(_01427_));
 sky130_fd_sc_hd__or2_1 _20590_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_03458_));
 sky130_fd_sc_hd__a32o_1 _20591_ (.A1(_07679_),
    .A2(_02830_),
    .A3(_03458_),
    .B1(_07855_),
    .B2(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_01428_));
 sky130_fd_sc_hd__a21bo_1 _20592_ (.A1(_02829_),
    .A2(_02831_),
    .B1_N(_02830_),
    .X(_03459_));
 sky130_fd_sc_hd__a32o_1 _20593_ (.A1(_07679_),
    .A2(_02832_),
    .A3(_03459_),
    .B1(_07855_),
    .B2(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_01429_));
 sky130_fd_sc_hd__and2b_1 _20594_ (.A_N(_02828_),
    .B(_02834_),
    .X(_03460_));
 sky130_fd_sc_hd__xnor2_1 _20595_ (.A(_02833_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a22o_1 _20596_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_03443_),
    .B1(_07756_),
    .B2(_03461_),
    .X(_01430_));
 sky130_fd_sc_hd__a21oi_1 _20597_ (.A1(_02827_),
    .A2(_02836_),
    .B1(_02835_),
    .Y(_03462_));
 sky130_fd_sc_hd__a31o_1 _20598_ (.A1(_02827_),
    .A2(_02836_),
    .A3(_02835_),
    .B1(_07830_),
    .X(_03463_));
 sky130_fd_sc_hd__a2bb2o_1 _20599_ (.A1_N(_03462_),
    .A2_N(_03463_),
    .B1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B2(_09762_),
    .X(_01431_));
 sky130_fd_sc_hd__nor2_1 _20600_ (.A(\gpout2.clk_div[0] ),
    .B(net60),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _20601_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .Y(_03464_));
 sky130_fd_sc_hd__or2_1 _20602_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .X(_03465_));
 sky130_fd_sc_hd__and3_1 _20603_ (.A(_02721_),
    .B(_03464_),
    .C(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _20604_ (.A(_03466_),
    .X(_01433_));
 sky130_fd_sc_hd__nor2_1 _20605_ (.A(\gpout3.clk_div[0] ),
    .B(net60),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_1 _20606_ (.A(\gpout3.clk_div[1] ),
    .B(\gpout3.clk_div[0] ),
    .Y(_03467_));
 sky130_fd_sc_hd__or2_1 _20607_ (.A(\gpout3.clk_div[1] ),
    .B(\gpout3.clk_div[0] ),
    .X(_03468_));
 sky130_fd_sc_hd__and3_1 _20608_ (.A(_02721_),
    .B(_03467_),
    .C(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _20609_ (.A(_03469_),
    .X(_01435_));
 sky130_fd_sc_hd__nor2_1 _20610_ (.A(\gpout4.clk_div[0] ),
    .B(net60),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_1 _20611_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .Y(_03470_));
 sky130_fd_sc_hd__or2_1 _20612_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .X(_03471_));
 sky130_fd_sc_hd__and3_1 _20613_ (.A(_02721_),
    .B(_03470_),
    .C(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _20614_ (.A(_03472_),
    .X(_01437_));
 sky130_fd_sc_hd__dfxtp_1 _20615_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00011_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20616_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00012_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20617_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00401_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_1 _20618_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00402_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_1 _20619_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00403_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_2 _20620_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00404_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_2 _20621_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00405_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20622_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20623_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00407_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_2 _20624_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00408_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_2 _20625_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00409_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _20626_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00410_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_2 _20627_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00411_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20628_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20629_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20630_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20631_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20632_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20633_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20634_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.mapY[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20635_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.stepDistY[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20636_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20637_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20638_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20639_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20640_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20641_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20642_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20643_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20644_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20645_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20646_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20647_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20648_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20649_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20650_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20651_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20652_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20653_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20654_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20655_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20656_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20657_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20658_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistY[11] ));
 sky130_fd_sc_hd__dfxtp_4 _20659_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.visualWallDist[-12] ));
 sky130_fd_sc_hd__dfxtp_4 _20660_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _20661_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _20662_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20663_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20664_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20665_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20666_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20667_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20668_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20669_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20670_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20671_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20672_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20673_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00457_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20674_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00458_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20675_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00459_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20676_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00460_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20677_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00461_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _20678_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00462_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20679_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00463_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_4 _20680_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00464_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_4 _20681_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00465_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20682_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00466_),
    .Q(\rbzero.wall_tracer.visualWallDist[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20683_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00467_),
    .Q(\rbzero.wall_tracer.stepDistX[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20684_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00468_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20685_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00469_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20686_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00470_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20687_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00471_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20688_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00472_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20689_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00473_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20690_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00474_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20691_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00475_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20692_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00476_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20693_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00477_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20694_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00478_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20695_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00479_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20696_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00480_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20697_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00481_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20698_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00482_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20699_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00483_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20700_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00484_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20701_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00485_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20702_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00486_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20703_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00487_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20704_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00488_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20705_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00489_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20706_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00490_),
    .Q(\rbzero.wall_tracer.stepDistX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20707_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00013_),
    .Q(\rbzero.wall_tracer.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20708_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00015_),
    .Q(\rbzero.wall_tracer.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20709_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20710_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20711_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00002_),
    .Q(\rbzero.wall_tracer.state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20712_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00003_),
    .Q(\rbzero.wall_tracer.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20713_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00004_),
    .Q(\rbzero.wall_tracer.state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20714_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00005_),
    .Q(\rbzero.wall_tracer.state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20715_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00016_),
    .Q(\rbzero.wall_tracer.state[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20716_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00006_),
    .Q(\rbzero.wall_tracer.state[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20717_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00007_),
    .Q(\rbzero.wall_tracer.state[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20718_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00008_),
    .Q(\rbzero.wall_tracer.state[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20719_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00009_),
    .Q(\rbzero.wall_tracer.state[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20720_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00010_),
    .Q(\rbzero.wall_tracer.state[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20721_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00014_),
    .Q(\rbzero.wall_tracer.state[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20722_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00491_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20723_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00492_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20724_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00493_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20725_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00494_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20726_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00495_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20727_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00496_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20728_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00497_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20729_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00498_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20730_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00499_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20731_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00500_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20732_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00501_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20733_ (.CLK(clknet_3_5_0_i_clk),
    .D(_00502_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20734_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00503_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20735_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00504_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20736_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00505_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20737_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00506_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20738_ (.CLK(clknet_3_5_0_i_clk),
    .D(_00507_),
    .Q(\rbzero.wall_tracer.rayAddendX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20739_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00508_),
    .Q(\rbzero.wall_tracer.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20740_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00509_),
    .Q(\rbzero.wall_tracer.wall[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20741_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00510_),
    .Q(\rbzero.wall_tracer.side ));
 sky130_fd_sc_hd__dfxtp_1 _20742_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00511_),
    .Q(\rbzero.wall_tracer.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20743_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00512_),
    .Q(\rbzero.wall_tracer.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20744_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00513_),
    .Q(\rbzero.wall_tracer.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20745_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00514_),
    .Q(\rbzero.wall_tracer.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20746_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00515_),
    .Q(\rbzero.wall_tracer.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20747_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00516_),
    .Q(\rbzero.wall_tracer.texu[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20748_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00517_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20749_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00518_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20750_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00519_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20751_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00520_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20752_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00521_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20753_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00522_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20754_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00523_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20755_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00524_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20756_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00525_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20757_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00526_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20758_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00527_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_2 _20759_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00528_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20760_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00529_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20761_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00530_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20762_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00531_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20763_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00532_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20764_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00533_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20765_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00534_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20766_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00535_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20767_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00536_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20768_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00537_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20769_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00538_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20770_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00539_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20771_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00540_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20772_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00541_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20773_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00542_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20774_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00543_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20775_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00544_),
    .Q(\rbzero.row_render.texu[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20776_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00545_),
    .Q(\rbzero.traced_texa[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20777_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00546_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20778_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00547_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20779_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00548_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20780_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00549_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20781_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00550_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20782_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00551_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20783_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00552_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20784_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00553_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20785_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00554_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20786_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00555_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20787_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00556_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20788_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00557_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20789_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00558_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20790_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00559_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20791_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00560_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20792_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00561_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20793_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00562_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20794_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00563_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20795_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00564_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20796_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00565_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20797_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00566_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20798_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00567_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20799_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00568_),
    .Q(\rbzero.traced_texa[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20800_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00569_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20801_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00570_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20802_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20803_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00572_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20804_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00573_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20805_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00574_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20806_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00575_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20807_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00576_),
    .Q(\rbzero.wall_tracer.mapX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20808_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00577_),
    .Q(\rbzero.wall_tracer.trackDistX[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20809_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00578_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20810_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00579_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20811_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00580_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20812_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00581_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20813_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00582_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20814_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00583_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20815_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00584_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20816_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00585_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20817_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00586_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20818_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00587_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20819_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00588_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20820_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00589_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20821_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00590_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20822_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00591_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20823_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00592_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20824_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00593_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20825_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00594_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20826_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00595_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20827_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00596_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20828_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00597_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20829_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00598_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20830_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00599_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20831_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00600_),
    .Q(\rbzero.wall_tracer.trackDistX[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20832_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00601_),
    .Q(\rbzero.wall_tracer.trackDistY[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _20833_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00602_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20834_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00603_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20835_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00604_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20836_ (.CLK(clknet_opt_10_1_i_clk),
    .D(_00605_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20837_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00606_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20838_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00607_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20839_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00608_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20840_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00609_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20841_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00610_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20842_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00611_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20843_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00612_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20844_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00613_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20845_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00614_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20846_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00615_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20847_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00616_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20848_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00617_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20849_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00618_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20850_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00619_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20851_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00620_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20852_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00621_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20853_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00622_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20854_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00623_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20855_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00624_),
    .Q(\rbzero.wall_tracer.trackDistY[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20856_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00625_),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _20857_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00626_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20858_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00627_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20859_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00628_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20860_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00629_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20861_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00630_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20862_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00631_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20863_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00632_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20864_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00633_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20865_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00634_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20866_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00635_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20867_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00636_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20868_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00637_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20869_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00638_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20870_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00639_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20871_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00640_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20872_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00641_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20873_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00642_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20874_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00643_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20875_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00644_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20876_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00645_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20877_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00646_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20878_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00647_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20879_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00648_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20880_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00649_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20881_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00650_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20882_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00651_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20883_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00652_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20884_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00653_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20885_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00654_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20886_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00655_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20887_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00656_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20888_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00657_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20889_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00658_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20890_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00659_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20891_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00660_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20892_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00661_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20893_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00662_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20894_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00663_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20895_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00664_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20896_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00665_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20897_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00666_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20898_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00667_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20899_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00668_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20900_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00669_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20901_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00670_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20902_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00671_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20903_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00672_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20904_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00673_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20905_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00674_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20906_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00675_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20907_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00676_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20908_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00677_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20909_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00678_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20910_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00679_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20911_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00680_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20912_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00681_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _20913_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00682_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20914_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00683_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20915_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00684_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20916_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00685_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20917_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00686_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20918_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00687_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00688_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20920_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00689_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00690_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20922_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00691_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20923_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00692_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20924_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00693_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00694_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20926_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00695_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00696_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20928_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00697_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _20929_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00698_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00699_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00700_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00701_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _20933_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00702_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00703_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _20935_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00704_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00705_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00706_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_2 _20938_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00707_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20939_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00708_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20940_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00709_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20941_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00710_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20942_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00711_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20943_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00712_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20944_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00713_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20945_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00714_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20946_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00715_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00716_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20948_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00717_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00718_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20950_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00719_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20951_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00720_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20952_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00721_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20953_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00722_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20954_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00723_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _20955_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00724_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20956_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00725_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20957_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00726_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20958_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00727_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20959_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00728_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20960_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00729_),
    .Q(\rbzero.otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20961_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00730_),
    .Q(\rbzero.otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20962_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00731_),
    .Q(\rbzero.otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20963_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00732_),
    .Q(\rbzero.otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20964_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00733_),
    .Q(\rbzero.otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20965_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00734_),
    .Q(\rbzero.othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20966_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00735_),
    .Q(\rbzero.othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20967_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00736_),
    .Q(\rbzero.othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00737_),
    .Q(\rbzero.othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00738_),
    .Q(\rbzero.othery[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20970_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00739_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00740_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00741_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00742_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00743_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00744_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00745_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00746_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00747_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00748_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00749_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00750_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00751_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00752_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20984_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00753_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00754_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00755_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00756_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00757_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00758_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00759_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00760_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20992_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00761_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20993_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00762_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20994_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00763_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00764_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _20996_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00765_),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20997_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00766_),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20998_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00767_),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20999_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00768_),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00769_),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21001_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00770_),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00771_),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _21003_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00772_),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00773_),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21005_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00774_),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00775_),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21007_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00776_),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00777_),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21009_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00778_),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _21010_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00779_),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21011_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00780_),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21012_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00781_),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21013_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00782_),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21014_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00783_),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21015_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00784_),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00785_),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00786_),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21018_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00787_),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00788_),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21020_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00789_),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00790_),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21022_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00791_),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00792_),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21024_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00793_),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21025_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00794_),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00795_),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21027_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00796_),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00797_),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21029_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00798_),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00799_),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21031_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00800_),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21032_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00801_),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00802_),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00803_),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00804_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00805_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21037_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00806_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00807_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21039_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00808_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00809_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00810_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00811_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21043_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00812_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00813_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00814_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21046_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00815_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21047_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00816_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00817_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00818_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21050_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00819_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00820_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21052_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00821_),
    .Q(\rbzero.wall_tracer.rayAddendY[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21053_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00822_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21054_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00823_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00824_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00825_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00826_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00827_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00828_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21060_ (.CLK(net150),
    .D(_00829_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(net151),
    .D(_00830_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(net152),
    .D(_00831_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(net153),
    .D(_00832_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(net154),
    .D(_00833_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(net155),
    .D(_00834_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(net156),
    .D(_00835_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(net157),
    .D(_00836_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(net158),
    .D(_00837_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(net159),
    .D(_00838_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(net160),
    .D(_00839_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(net161),
    .D(_00840_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(net162),
    .D(_00841_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(net163),
    .D(_00842_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(net164),
    .D(_00843_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(net165),
    .D(_00844_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(net166),
    .D(_00845_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(net167),
    .D(_00846_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(net168),
    .D(_00847_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(net169),
    .D(_00848_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(net170),
    .D(_00849_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(net171),
    .D(_00850_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(net172),
    .D(_00851_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(net173),
    .D(_00852_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(net174),
    .D(_00853_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(net175),
    .D(_00854_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(net176),
    .D(_00855_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(net177),
    .D(_00856_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(net178),
    .D(_00857_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(net179),
    .D(_00858_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(net180),
    .D(_00859_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(net181),
    .D(_00860_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21092_ (.CLK(net182),
    .D(_00861_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(net183),
    .D(_00862_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(net184),
    .D(_00863_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(net185),
    .D(_00864_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(net186),
    .D(_00865_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(net187),
    .D(_00866_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21098_ (.CLK(net188),
    .D(_00867_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21099_ (.CLK(net189),
    .D(_00868_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(net190),
    .D(_00869_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21101_ (.CLK(net191),
    .D(_00870_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21102_ (.CLK(net192),
    .D(_00871_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(net193),
    .D(_00872_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21104_ (.CLK(net194),
    .D(_00873_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(net195),
    .D(_00874_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(net196),
    .D(_00875_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21107_ (.CLK(net197),
    .D(_00876_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(net198),
    .D(_00877_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(net199),
    .D(_00878_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(net200),
    .D(_00879_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21111_ (.CLK(net201),
    .D(_00880_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21112_ (.CLK(net202),
    .D(_00881_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21113_ (.CLK(net203),
    .D(_00882_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(net204),
    .D(_00883_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21115_ (.CLK(net205),
    .D(_00884_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21116_ (.CLK(net206),
    .D(_00885_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21117_ (.CLK(net207),
    .D(_00886_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(net208),
    .D(_00887_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21119_ (.CLK(net209),
    .D(_00888_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21120_ (.CLK(net210),
    .D(_00889_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(net211),
    .D(_00890_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(net212),
    .D(_00891_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(net213),
    .D(_00892_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00893_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00894_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00895_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00896_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00897_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21129_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00898_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21130_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00899_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00900_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00901_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00902_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00903_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00904_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21136_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00905_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00906_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00907_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21139_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00908_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21140_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00909_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21141_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00910_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21142_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00911_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21143_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00912_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21144_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00913_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21145_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00914_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21146_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00915_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21147_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00916_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21148_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00917_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21149_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00918_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21150_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00919_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21151_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00920_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21152_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00921_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21153_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00922_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00923_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21155_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00924_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21156_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00925_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00926_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21158_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00927_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21159_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00928_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00929_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00930_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21162_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00931_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21163_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00932_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00933_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00934_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21166_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00935_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00936_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00937_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00938_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00939_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00940_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00941_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00942_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00943_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00944_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21176_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00945_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00946_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00947_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00948_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00949_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00950_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00951_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00952_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00953_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00954_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00955_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00956_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00957_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00958_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00959_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00960_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00961_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00962_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00963_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00964_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00965_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00966_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00967_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00968_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00969_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00970_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00971_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00972_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00973_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21205_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00974_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21206_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00975_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00976_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00977_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21209_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00978_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00979_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00980_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21212_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00981_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00982_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21214_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00983_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21215_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00984_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21216_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00985_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21217_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00986_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00987_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00988_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21220_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00989_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21221_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00990_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00991_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00992_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00993_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21225_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00994_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21226_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00995_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21227_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00996_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00997_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21229_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00998_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21230_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00999_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21231_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01000_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21232_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01001_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21233_ (.CLK(clknet_leaf_18_i_clk),
    .D(_01002_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21234_ (.CLK(clknet_leaf_18_i_clk),
    .D(_01003_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01004_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01005_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01006_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01007_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21239_ (.CLK(clknet_leaf_68_i_clk),
    .D(_01008_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21240_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01009_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21241_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01010_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01011_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21243_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01012_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01013_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21245_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01014_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01015_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21247_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01016_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21248_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01017_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21249_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01018_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21250_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01019_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21251_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01020_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21252_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01021_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21253_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01022_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21254_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01023_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21255_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01024_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21256_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01025_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21257_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01026_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21258_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01027_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_4 _21259_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01028_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21260_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01029_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_4 _21261_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01030_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_4 _21262_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01031_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01032_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _21264_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01033_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01034_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01035_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21267_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01036_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21268_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01037_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21269_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01038_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_4 _21270_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01039_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21271_ (.CLK(clknet_leaf_5_i_clk),
    .D(_01040_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21272_ (.CLK(clknet_leaf_5_i_clk),
    .D(_01041_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21273_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01042_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01043_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _21275_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01044_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _21276_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01045_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_4 _21277_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01046_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21278_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01047_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01048_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_2 _21280_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01049_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01050_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01051_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01052_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01053_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21285_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01054_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_4 _21286_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01055_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_4 _21287_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01056_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01057_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01058_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01059_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01060_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_3_i_clk),
    .D(_01061_),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(net214),
    .D(_01062_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(net215),
    .D(_01063_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(net216),
    .D(_01064_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(net217),
    .D(_01065_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(net218),
    .D(_01066_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(net219),
    .D(_01067_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(net220),
    .D(_01068_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(net221),
    .D(_01069_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(net222),
    .D(_01070_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(net223),
    .D(_01071_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(net224),
    .D(_01072_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(net225),
    .D(_01073_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(net226),
    .D(_01074_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(net227),
    .D(_01075_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(net228),
    .D(_01076_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(net229),
    .D(_01077_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(net230),
    .D(_01078_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(net231),
    .D(_01079_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(net232),
    .D(_01080_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(net233),
    .D(_01081_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(net234),
    .D(_01082_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(net235),
    .D(_01083_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(net236),
    .D(_01084_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(net237),
    .D(_01085_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(net238),
    .D(_01086_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(net239),
    .D(_01087_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(net240),
    .D(_01088_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(net241),
    .D(_01089_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(net242),
    .D(_01090_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(net243),
    .D(_01091_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(net244),
    .D(_01092_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(net245),
    .D(_01093_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(net246),
    .D(_01094_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(net247),
    .D(_01095_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(net248),
    .D(_01096_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(net249),
    .D(_01097_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(net250),
    .D(_01098_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(net251),
    .D(_01099_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(net252),
    .D(_01100_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(net253),
    .D(_01101_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(net254),
    .D(_01102_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(net255),
    .D(_01103_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(net256),
    .D(_01104_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(net257),
    .D(_01105_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(net258),
    .D(_01106_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(net259),
    .D(_01107_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(net260),
    .D(_01108_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(net261),
    .D(_01109_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(net262),
    .D(_01110_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(net263),
    .D(_01111_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(net264),
    .D(_01112_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(net265),
    .D(_01113_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(net266),
    .D(_01114_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(net267),
    .D(_01115_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(net268),
    .D(_01116_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(net269),
    .D(_01117_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(net270),
    .D(_01118_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(net271),
    .D(_01119_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(net272),
    .D(_01120_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(net273),
    .D(_01121_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(net274),
    .D(_01122_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(net275),
    .D(_01123_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(net276),
    .D(_01124_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(net277),
    .D(_01125_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(net278),
    .D(_01126_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(net279),
    .D(_01127_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(net280),
    .D(_01128_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(net281),
    .D(_01129_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(net282),
    .D(_01130_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(net283),
    .D(_01131_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(net284),
    .D(_01132_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(net285),
    .D(_01133_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(net286),
    .D(_01134_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(net287),
    .D(_01135_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(net288),
    .D(_01136_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(net289),
    .D(_01137_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(net290),
    .D(_01138_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(net291),
    .D(_01139_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(net292),
    .D(_01140_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(net293),
    .D(_01141_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(net294),
    .D(_01142_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(net295),
    .D(_01143_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(net296),
    .D(_01144_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(net297),
    .D(_01145_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(net298),
    .D(_01146_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(net299),
    .D(_01147_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(net300),
    .D(_01148_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(net301),
    .D(_01149_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(net302),
    .D(_01150_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(net303),
    .D(_01151_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(net304),
    .D(_01152_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(net305),
    .D(_01153_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(net306),
    .D(_01154_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(net307),
    .D(_01155_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(net308),
    .D(_01156_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(net309),
    .D(_01157_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(net310),
    .D(_01158_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(net311),
    .D(_01159_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(net312),
    .D(_01160_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(net313),
    .D(_01161_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(net314),
    .D(_01162_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(net315),
    .D(_01163_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(net316),
    .D(_01164_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(net317),
    .D(_01165_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(net318),
    .D(_01166_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(net319),
    .D(_01167_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(net320),
    .D(_01168_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(net321),
    .D(_01169_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(net322),
    .D(_01170_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(net323),
    .D(_01171_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(net324),
    .D(_01172_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(net325),
    .D(_01173_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(net326),
    .D(_01174_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(net327),
    .D(_01175_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(net328),
    .D(_01176_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(net329),
    .D(_01177_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(net330),
    .D(_01178_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(net331),
    .D(_01179_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(net332),
    .D(_01180_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(net333),
    .D(_01181_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(net334),
    .D(_01182_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(net335),
    .D(_01183_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(net336),
    .D(_01184_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(net337),
    .D(_01185_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(net338),
    .D(_01186_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(net339),
    .D(_01187_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21419_ (.CLK(net340),
    .D(_01188_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(net341),
    .D(_01189_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(net342),
    .D(_01190_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(net343),
    .D(_01191_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(net344),
    .D(_01192_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(net345),
    .D(_01193_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(net346),
    .D(_01194_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(net347),
    .D(_01195_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(net348),
    .D(_01196_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(net349),
    .D(_01197_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(net350),
    .D(_01198_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(net351),
    .D(_01199_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(net352),
    .D(_01200_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(net353),
    .D(_01201_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21433_ (.CLK(net354),
    .D(_01202_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21434_ (.CLK(net355),
    .D(_01203_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(net356),
    .D(_01204_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(net357),
    .D(_01205_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(net358),
    .D(_01206_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(net359),
    .D(_01207_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(net360),
    .D(_01208_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(net361),
    .D(_01209_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21441_ (.CLK(net362),
    .D(_01210_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(net363),
    .D(_01211_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(net364),
    .D(_01212_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(net365),
    .D(_01213_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(net366),
    .D(_01214_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(net367),
    .D(_01215_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(net368),
    .D(_01216_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(net369),
    .D(_01217_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(net370),
    .D(_01218_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(net371),
    .D(_01219_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(net372),
    .D(_01220_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(net373),
    .D(_01221_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(net374),
    .D(_01222_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(net375),
    .D(_01223_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(net376),
    .D(_01224_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(net377),
    .D(_01225_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(net378),
    .D(_01226_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(net379),
    .D(_01227_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(net380),
    .D(_01228_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(net381),
    .D(_01229_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(net382),
    .D(_01230_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(net383),
    .D(_01231_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(net384),
    .D(_01232_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(net385),
    .D(_01233_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(net386),
    .D(_01234_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(net387),
    .D(_01235_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(net388),
    .D(_01236_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(net389),
    .D(_01237_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(net390),
    .D(_01238_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(net391),
    .D(_01239_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(net392),
    .D(_01240_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(net393),
    .D(_01241_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(net394),
    .D(_01242_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(net395),
    .D(_01243_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(net396),
    .D(_01244_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(net397),
    .D(_01245_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(net398),
    .D(_01246_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(net399),
    .D(_01247_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(net400),
    .D(_01248_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(net401),
    .D(_01249_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(net402),
    .D(_01250_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(net403),
    .D(_01251_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(net404),
    .D(_01252_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(net405),
    .D(_01253_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(net406),
    .D(_01254_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21486_ (.CLK(net407),
    .D(_01255_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(net408),
    .D(_01256_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(net409),
    .D(_01257_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(net410),
    .D(_01258_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(net411),
    .D(_01259_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21491_ (.CLK(net412),
    .D(_01260_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(net413),
    .D(_01261_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(net414),
    .D(_01262_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(net415),
    .D(_01263_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(net416),
    .D(_01264_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(net417),
    .D(_01265_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(net418),
    .D(_01266_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(net419),
    .D(_01267_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(net420),
    .D(_01268_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(net421),
    .D(_01269_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(net422),
    .D(_01270_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21502_ (.CLK(net423),
    .D(_01271_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(net424),
    .D(_01272_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(net425),
    .D(_01273_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(net426),
    .D(_01274_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(net427),
    .D(_01275_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(net428),
    .D(_01276_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(net429),
    .D(_01277_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(net430),
    .D(_01278_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(net431),
    .D(_01279_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(net432),
    .D(_01280_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(net433),
    .D(_01281_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(net434),
    .D(_01282_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(net435),
    .D(_01283_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(net436),
    .D(_01284_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(net437),
    .D(_01285_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(net438),
    .D(_01286_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(net439),
    .D(_01287_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(net440),
    .D(_01288_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(net441),
    .D(_01289_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(net442),
    .D(_01290_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(net443),
    .D(_01291_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(net444),
    .D(_01292_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(net445),
    .D(_01293_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(net446),
    .D(_01294_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(net447),
    .D(_01295_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(net448),
    .D(_01296_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(net449),
    .D(_01297_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(net450),
    .D(_01298_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(net451),
    .D(_01299_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(net452),
    .D(_01300_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(net453),
    .D(_01301_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(net454),
    .D(_01302_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(net455),
    .D(_01303_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(net456),
    .D(_01304_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(net457),
    .D(_01305_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(net458),
    .D(_01306_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(net459),
    .D(_01307_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(net460),
    .D(_01308_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(net461),
    .D(_01309_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(net462),
    .D(_01310_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(net463),
    .D(_01311_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(net464),
    .D(_01312_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(net465),
    .D(_01313_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(net466),
    .D(_01314_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(net467),
    .D(_01315_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(net468),
    .D(_01316_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(net469),
    .D(_01317_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(net470),
    .D(_01318_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(net471),
    .D(_01319_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(net472),
    .D(_01320_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(net473),
    .D(_01321_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(net474),
    .D(_01322_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(net475),
    .D(_01323_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(net476),
    .D(_01324_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(net477),
    .D(_01325_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21557_ (.CLK(net478),
    .D(_01326_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(net479),
    .D(_01327_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21559_ (.CLK(net480),
    .D(_01328_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(net481),
    .D(_01329_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(net482),
    .D(_01330_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(net483),
    .D(_01331_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(net484),
    .D(_01332_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(net485),
    .D(_01333_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(net486),
    .D(_01334_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(net487),
    .D(_01335_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(net488),
    .D(_01336_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(net489),
    .D(_01337_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(net490),
    .D(_01338_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(net491),
    .D(_01339_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(net492),
    .D(_01340_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(net493),
    .D(_01341_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(net494),
    .D(_01342_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(net495),
    .D(_01343_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(net496),
    .D(_01344_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(net497),
    .D(_01345_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(net498),
    .D(_01346_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(net499),
    .D(_01347_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(net500),
    .D(_01348_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(net501),
    .D(_01349_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(net502),
    .D(_01350_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21582_ (.CLK(net503),
    .D(_01351_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(net504),
    .D(_01352_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(net505),
    .D(_01353_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(net506),
    .D(_01354_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(net507),
    .D(_01355_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(net508),
    .D(_01356_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(net509),
    .D(_01357_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(net130),
    .D(_01358_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(net131),
    .D(_01359_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(net132),
    .D(_01360_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(net133),
    .D(_01361_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21593_ (.CLK(net134),
    .D(_01362_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(net135),
    .D(_01363_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(net136),
    .D(_01364_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(net137),
    .D(_01365_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(net138),
    .D(_01366_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(net139),
    .D(_01367_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(net140),
    .D(_01368_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21600_ (.CLK(net141),
    .D(_01369_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(net142),
    .D(_01370_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(net143),
    .D(_01371_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21603_ (.CLK(net144),
    .D(_01372_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(net145),
    .D(_01373_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21605_ (.CLK(net146),
    .D(_01374_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(net147),
    .D(_01375_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(net148),
    .D(_01376_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(net149),
    .D(_01377_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(net126),
    .D(_01378_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(net127),
    .D(_01379_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(net128),
    .D(_01380_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(net129),
    .D(_01381_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01382_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21614_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01383_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01384_),
    .Q(\rbzero.texV[-12] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01385_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01386_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01387_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01388_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01389_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01390_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01391_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01392_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01393_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01394_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01395_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01396_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01397_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01398_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01399_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21631_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01400_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21632_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01401_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01402_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21634_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01403_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21635_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01404_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21636_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01405_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01406_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21638_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01407_),
    .Q(\rbzero.texV[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01408_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01409_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21641_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01410_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01411_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01412_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01413_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21645_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01414_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21646_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01415_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01416_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01417_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21649_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01418_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01419_),
    .Q(\rbzero.traced_texVinit[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21651_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01420_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01421_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01422_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01423_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01424_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01425_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01426_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01427_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01428_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01429_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01430_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01431_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01432_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01433_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01434_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01435_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01436_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01437_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.HI(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.HI(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.HI(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.HI(net110));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.HI(net121));
 sky130_fd_sc_hd__inv_2 _12063__1 (.A(clknet_1_1__leaf__04835_),
    .Y(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.HI(net106));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(i_debug_vec_overlay),
    .X(net1));
 sky130_fd_sc_hd__buf_8 input2 (.A(i_gpout0_sel[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_8 input3 (.A(i_gpout0_sel[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_8 input4 (.A(i_gpout0_sel[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_8 input5 (.A(i_gpout0_sel[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_8 input6 (.A(i_gpout0_sel[4]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(i_gpout0_sel[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 input8 (.A(i_gpout1_sel[0]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout1_sel[1]),
    .X(net9));
 sky130_fd_sc_hd__buf_8 input10 (.A(i_gpout1_sel[2]),
    .X(net10));
 sky130_fd_sc_hd__buf_8 input11 (.A(i_gpout1_sel[3]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(i_gpout1_sel[4]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(i_gpout1_sel[5]),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input14 (.A(i_gpout2_sel[0]),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(i_gpout2_sel[1]),
    .X(net15));
 sky130_fd_sc_hd__buf_8 input16 (.A(i_gpout2_sel[2]),
    .X(net16));
 sky130_fd_sc_hd__buf_8 input17 (.A(i_gpout2_sel[3]),
    .X(net17));
 sky130_fd_sc_hd__buf_8 input18 (.A(i_gpout2_sel[4]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(i_gpout2_sel[5]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input20 (.A(i_gpout3_sel[0]),
    .X(net20));
 sky130_fd_sc_hd__buf_6 input21 (.A(i_gpout3_sel[1]),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input22 (.A(i_gpout3_sel[2]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(i_gpout3_sel[3]),
    .X(net23));
 sky130_fd_sc_hd__buf_6 input24 (.A(i_gpout3_sel[4]),
    .X(net24));
 sky130_fd_sc_hd__buf_6 input25 (.A(i_gpout3_sel[5]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(i_gpout4_sel[0]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(i_gpout4_sel[1]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 input28 (.A(i_gpout4_sel[2]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(i_gpout4_sel[3]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input30 (.A(i_gpout4_sel[4]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(i_gpout4_sel[5]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(i_gpout5_sel[0]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(i_gpout5_sel[1]),
    .X(net33));
 sky130_fd_sc_hd__buf_6 input34 (.A(i_gpout5_sel[2]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(i_gpout5_sel[3]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(i_gpout5_sel[4]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(i_gpout5_sel[5]),
    .X(net37));
 sky130_fd_sc_hd__buf_8 input38 (.A(i_mode[0]),
    .X(net38));
 sky130_fd_sc_hd__buf_8 input39 (.A(i_mode[1]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input40 (.A(i_mode[2]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_16 input41 (.A(i_reg_csb),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_16 input42 (.A(i_reg_mosi),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(i_reg_sclk),
    .X(net43));
 sky130_fd_sc_hd__buf_6 input44 (.A(i_reset_lock_a),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(i_reset_lock_b),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(i_tex_in[0]),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(i_tex_in[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_tex_in[2]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(i_tex_in[3]),
    .X(net49));
 sky130_fd_sc_hd__buf_8 input50 (.A(i_vec_csb),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(i_vec_mosi),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(i_vec_sclk),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net510),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(o_hsync));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(o_reset));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(o_tex_csb));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(o_tex_out0));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net122),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(o_vsync));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_72 (.LO(net72));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_1_1__leaf__04835_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 net99_3 (.A(clknet_1_1__leaf__04835_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 net99_4 (.A(clknet_1_1__leaf__04835_),
    .Y(net125));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_opt_4_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_opt_6_1_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_opt_7_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_opt_8_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_opt_9_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_opt_12_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_opt_13_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_opt_11_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_opt_2_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_opt_3_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_opt_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_opt_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_opt_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_1_i_clk (.A(clknet_opt_6_0_i_clk),
    .X(clknet_opt_6_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_9_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_opt_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_1_i_clk (.A(clknet_opt_10_0_i_clk),
    .X(clknet_opt_10_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_11_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_opt_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_12_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_opt_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_13_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_opt_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04835_ (.A(_04835_),
    .X(clknet_0__04835_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04835_ (.A(clknet_0__04835_),
    .X(clknet_1_0__leaf__04835_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04835_ (.A(clknet_0__04835_),
    .X(clknet_1_1__leaf__04835_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03321_ (.A(_03321_),
    .X(clknet_0__03321_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03321_ (.A(clknet_0__03321_),
    .X(clknet_1_0__leaf__03321_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03321_ (.A(clknet_0__03321_),
    .X(clknet_1_1__leaf__03321_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03320_ (.A(_03320_),
    .X(clknet_0__03320_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03320_ (.A(clknet_0__03320_),
    .X(clknet_1_0__leaf__03320_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03320_ (.A(clknet_0__03320_),
    .X(clknet_1_1__leaf__03320_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03309_ (.A(_03309_),
    .X(clknet_0__03309_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03309_ (.A(clknet_0__03309_),
    .X(clknet_1_0__leaf__03309_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03309_ (.A(clknet_0__03309_),
    .X(clknet_1_1__leaf__03309_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03319_ (.A(_03319_),
    .X(clknet_0__03319_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03319_ (.A(clknet_0__03319_),
    .X(clknet_1_0__leaf__03319_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03319_ (.A(clknet_0__03319_),
    .X(clknet_1_1__leaf__03319_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03318_ (.A(_03318_),
    .X(clknet_0__03318_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03318_ (.A(clknet_0__03318_),
    .X(clknet_1_0__leaf__03318_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03318_ (.A(clknet_0__03318_),
    .X(clknet_1_1__leaf__03318_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03317_ (.A(_03317_),
    .X(clknet_0__03317_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03317_ (.A(clknet_0__03317_),
    .X(clknet_1_0__leaf__03317_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03317_ (.A(clknet_0__03317_),
    .X(clknet_1_1__leaf__03317_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03316_ (.A(_03316_),
    .X(clknet_0__03316_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03316_ (.A(clknet_0__03316_),
    .X(clknet_1_0__leaf__03316_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03316_ (.A(clknet_0__03316_),
    .X(clknet_1_1__leaf__03316_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03315_ (.A(_03315_),
    .X(clknet_0__03315_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03315_ (.A(clknet_0__03315_),
    .X(clknet_1_0__leaf__03315_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03315_ (.A(clknet_0__03315_),
    .X(clknet_1_1__leaf__03315_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03314_ (.A(_03314_),
    .X(clknet_0__03314_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03314_ (.A(clknet_0__03314_),
    .X(clknet_1_0__leaf__03314_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03314_ (.A(clknet_0__03314_),
    .X(clknet_1_1__leaf__03314_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03313_ (.A(_03313_),
    .X(clknet_0__03313_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03313_ (.A(clknet_0__03313_),
    .X(clknet_1_0__leaf__03313_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03313_ (.A(clknet_0__03313_),
    .X(clknet_1_1__leaf__03313_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03312_ (.A(_03312_),
    .X(clknet_0__03312_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03312_ (.A(clknet_0__03312_),
    .X(clknet_1_0__leaf__03312_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03312_ (.A(clknet_0__03312_),
    .X(clknet_1_1__leaf__03312_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03311_ (.A(_03311_),
    .X(clknet_0__03311_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03311_ (.A(clknet_0__03311_),
    .X(clknet_1_0__leaf__03311_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03311_ (.A(clknet_0__03311_),
    .X(clknet_1_1__leaf__03311_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03310_ (.A(_03310_),
    .X(clknet_0__03310_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03310_ (.A(clknet_0__03310_),
    .X(clknet_1_0__leaf__03310_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03310_ (.A(clknet_0__03310_),
    .X(clknet_1_1__leaf__03310_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03298_ (.A(_03298_),
    .X(clknet_0__03298_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03298_ (.A(clknet_0__03298_),
    .X(clknet_1_0__leaf__03298_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03298_ (.A(clknet_0__03298_),
    .X(clknet_1_1__leaf__03298_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03308_ (.A(_03308_),
    .X(clknet_0__03308_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03308_ (.A(clknet_0__03308_),
    .X(clknet_1_0__leaf__03308_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03308_ (.A(clknet_0__03308_),
    .X(clknet_1_1__leaf__03308_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03307_ (.A(_03307_),
    .X(clknet_0__03307_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03307_ (.A(clknet_0__03307_),
    .X(clknet_1_0__leaf__03307_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03307_ (.A(clknet_0__03307_),
    .X(clknet_1_1__leaf__03307_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03306_ (.A(_03306_),
    .X(clknet_0__03306_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03306_ (.A(clknet_0__03306_),
    .X(clknet_1_0__leaf__03306_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03306_ (.A(clknet_0__03306_),
    .X(clknet_1_1__leaf__03306_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03305_ (.A(_03305_),
    .X(clknet_0__03305_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03305_ (.A(clknet_0__03305_),
    .X(clknet_1_0__leaf__03305_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03305_ (.A(clknet_0__03305_),
    .X(clknet_1_1__leaf__03305_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03304_ (.A(_03304_),
    .X(clknet_0__03304_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03304_ (.A(clknet_0__03304_),
    .X(clknet_1_0__leaf__03304_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03304_ (.A(clknet_0__03304_),
    .X(clknet_1_1__leaf__03304_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03303_ (.A(_03303_),
    .X(clknet_0__03303_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03303_ (.A(clknet_0__03303_),
    .X(clknet_1_0__leaf__03303_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03303_ (.A(clknet_0__03303_),
    .X(clknet_1_1__leaf__03303_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03302_ (.A(_03302_),
    .X(clknet_0__03302_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03302_ (.A(clknet_0__03302_),
    .X(clknet_1_0__leaf__03302_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03302_ (.A(clknet_0__03302_),
    .X(clknet_1_1__leaf__03302_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03301_ (.A(_03301_),
    .X(clknet_0__03301_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03301_ (.A(clknet_0__03301_),
    .X(clknet_1_0__leaf__03301_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03301_ (.A(clknet_0__03301_),
    .X(clknet_1_1__leaf__03301_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03300_ (.A(_03300_),
    .X(clknet_0__03300_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03300_ (.A(clknet_0__03300_),
    .X(clknet_1_0__leaf__03300_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03300_ (.A(clknet_0__03300_),
    .X(clknet_1_1__leaf__03300_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03299_ (.A(_03299_),
    .X(clknet_0__03299_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03299_ (.A(clknet_0__03299_),
    .X(clknet_1_0__leaf__03299_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03299_ (.A(clknet_0__03299_),
    .X(clknet_1_1__leaf__03299_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03044_ (.A(_03044_),
    .X(clknet_0__03044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03044_ (.A(clknet_0__03044_),
    .X(clknet_1_0__leaf__03044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03044_ (.A(clknet_0__03044_),
    .X(clknet_1_1__leaf__03044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03297_ (.A(_03297_),
    .X(clknet_0__03297_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03297_ (.A(clknet_0__03297_),
    .X(clknet_1_0__leaf__03297_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03297_ (.A(clknet_0__03297_),
    .X(clknet_1_1__leaf__03297_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03296_ (.A(_03296_),
    .X(clknet_0__03296_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03296_ (.A(clknet_0__03296_),
    .X(clknet_1_0__leaf__03296_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03296_ (.A(clknet_0__03296_),
    .X(clknet_1_1__leaf__03296_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03295_ (.A(_03295_),
    .X(clknet_0__03295_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03295_ (.A(clknet_0__03295_),
    .X(clknet_1_0__leaf__03295_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03295_ (.A(clknet_0__03295_),
    .X(clknet_1_1__leaf__03295_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03294_ (.A(_03294_),
    .X(clknet_0__03294_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03294_ (.A(clknet_0__03294_),
    .X(clknet_1_0__leaf__03294_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03294_ (.A(clknet_0__03294_),
    .X(clknet_1_1__leaf__03294_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03293_ (.A(_03293_),
    .X(clknet_0__03293_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03293_ (.A(clknet_0__03293_),
    .X(clknet_1_0__leaf__03293_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03293_ (.A(clknet_0__03293_),
    .X(clknet_1_1__leaf__03293_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03292_ (.A(_03292_),
    .X(clknet_0__03292_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03292_ (.A(clknet_0__03292_),
    .X(clknet_1_0__leaf__03292_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03292_ (.A(clknet_0__03292_),
    .X(clknet_1_1__leaf__03292_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03291_ (.A(_03291_),
    .X(clknet_0__03291_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03291_ (.A(clknet_0__03291_),
    .X(clknet_1_0__leaf__03291_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03291_ (.A(clknet_0__03291_),
    .X(clknet_1_1__leaf__03291_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03290_ (.A(_03290_),
    .X(clknet_0__03290_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03290_ (.A(clknet_0__03290_),
    .X(clknet_1_0__leaf__03290_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03290_ (.A(clknet_0__03290_),
    .X(clknet_1_1__leaf__03290_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03289_ (.A(_03289_),
    .X(clknet_0__03289_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03289_ (.A(clknet_0__03289_),
    .X(clknet_1_0__leaf__03289_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03289_ (.A(clknet_0__03289_),
    .X(clknet_1_1__leaf__03289_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03045_ (.A(_03045_),
    .X(clknet_0__03045_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03045_ (.A(clknet_0__03045_),
    .X(clknet_1_0__leaf__03045_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03045_ (.A(clknet_0__03045_),
    .X(clknet_1_1__leaf__03045_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03037_ (.A(_03037_),
    .X(clknet_0__03037_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03037_ (.A(clknet_0__03037_),
    .X(clknet_1_0__leaf__03037_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03037_ (.A(clknet_0__03037_),
    .X(clknet_1_1__leaf__03037_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03043_ (.A(_03043_),
    .X(clknet_0__03043_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03043_ (.A(clknet_0__03043_),
    .X(clknet_1_0__leaf__03043_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03043_ (.A(clknet_0__03043_),
    .X(clknet_1_1__leaf__03043_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03042_ (.A(_03042_),
    .X(clknet_0__03042_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03042_ (.A(clknet_0__03042_),
    .X(clknet_1_0__leaf__03042_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03042_ (.A(clknet_0__03042_),
    .X(clknet_1_1__leaf__03042_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03041_ (.A(_03041_),
    .X(clknet_0__03041_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03041_ (.A(clknet_0__03041_),
    .X(clknet_1_0__leaf__03041_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03041_ (.A(clknet_0__03041_),
    .X(clknet_1_1__leaf__03041_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03040_ (.A(_03040_),
    .X(clknet_0__03040_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03040_ (.A(clknet_0__03040_),
    .X(clknet_1_0__leaf__03040_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03040_ (.A(clknet_0__03040_),
    .X(clknet_1_1__leaf__03040_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03039_ (.A(_03039_),
    .X(clknet_0__03039_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03039_ (.A(clknet_0__03039_),
    .X(clknet_1_0__leaf__03039_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03039_ (.A(clknet_0__03039_),
    .X(clknet_1_1__leaf__03039_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03038_ (.A(_03038_),
    .X(clknet_0__03038_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03038_ (.A(clknet_0__03038_),
    .X(clknet_1_0__leaf__03038_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03038_ (.A(clknet_0__03038_),
    .X(clknet_1_1__leaf__03038_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rbzero.tex_r1[40] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rbzero.pov.ready_buffer[31] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\rbzero.wall_tracer.texu[3] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\rbzero.pov.spi_buffer[31] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\rbzero.pov.ready_buffer[29] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_05190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_05204_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_05533_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_05893_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_07514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_07524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_07524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_07530_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_07541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_08037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_08039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_08094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_08283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_09162_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_09350_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_09611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_09765_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_09781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_09807_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\rbzero.wall_tracer.visualWallDist[-12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_07536_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_07549_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_07916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_07939_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_08159_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_09859_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_10297_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net66));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_980 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1229 ();
 assign o_rgb[0] = net72;
 assign o_rgb[10] = net80;
 assign o_rgb[11] = net81;
 assign o_rgb[12] = net82;
 assign o_rgb[13] = net83;
 assign o_rgb[16] = net84;
 assign o_rgb[17] = net85;
 assign o_rgb[18] = net86;
 assign o_rgb[19] = net87;
 assign o_rgb[1] = net73;
 assign o_rgb[20] = net88;
 assign o_rgb[21] = net89;
 assign o_rgb[2] = net74;
 assign o_rgb[3] = net75;
 assign o_rgb[4] = net76;
 assign o_rgb[5] = net77;
 assign o_rgb[8] = net78;
 assign o_rgb[9] = net79;
 assign ones[0] = net106;
 assign ones[10] = net116;
 assign ones[11] = net117;
 assign ones[12] = net118;
 assign ones[13] = net119;
 assign ones[14] = net120;
 assign ones[15] = net121;
 assign ones[1] = net107;
 assign ones[2] = net108;
 assign ones[3] = net109;
 assign ones[4] = net110;
 assign ones[5] = net111;
 assign ones[6] = net112;
 assign ones[7] = net113;
 assign ones[8] = net114;
 assign ones[9] = net115;
 assign zeros[0] = net90;
 assign zeros[10] = net100;
 assign zeros[11] = net101;
 assign zeros[12] = net102;
 assign zeros[13] = net103;
 assign zeros[14] = net104;
 assign zeros[15] = net105;
 assign zeros[1] = net91;
 assign zeros[2] = net92;
 assign zeros[3] = net93;
 assign zeros[4] = net94;
 assign zeros[5] = net95;
 assign zeros[6] = net96;
 assign zeros[7] = net97;
 assign zeros[8] = net98;
 assign zeros[9] = net99;
endmodule


magic
tech sky130A
magscale 1 2
timestamp 1698657145
<< viali >>
rect 14473 43673 14507 43707
rect 14473 35989 14507 36023
rect 14473 27965 14507 27999
rect 14473 20349 14507 20383
rect 14473 12121 14507 12155
rect 14473 4437 14507 4471
<< metal1 >>
rect 1104 45722 14971 45744
rect 1104 45670 4376 45722
rect 4428 45670 4440 45722
rect 4492 45670 4504 45722
rect 4556 45670 4568 45722
rect 4620 45670 4632 45722
rect 4684 45670 7803 45722
rect 7855 45670 7867 45722
rect 7919 45670 7931 45722
rect 7983 45670 7995 45722
rect 8047 45670 8059 45722
rect 8111 45670 11230 45722
rect 11282 45670 11294 45722
rect 11346 45670 11358 45722
rect 11410 45670 11422 45722
rect 11474 45670 11486 45722
rect 11538 45670 14657 45722
rect 14709 45670 14721 45722
rect 14773 45670 14785 45722
rect 14837 45670 14849 45722
rect 14901 45670 14913 45722
rect 14965 45670 14971 45722
rect 1104 45648 14971 45670
rect 1104 45178 14812 45200
rect 1104 45126 2663 45178
rect 2715 45126 2727 45178
rect 2779 45126 2791 45178
rect 2843 45126 2855 45178
rect 2907 45126 2919 45178
rect 2971 45126 6090 45178
rect 6142 45126 6154 45178
rect 6206 45126 6218 45178
rect 6270 45126 6282 45178
rect 6334 45126 6346 45178
rect 6398 45126 9517 45178
rect 9569 45126 9581 45178
rect 9633 45126 9645 45178
rect 9697 45126 9709 45178
rect 9761 45126 9773 45178
rect 9825 45126 12944 45178
rect 12996 45126 13008 45178
rect 13060 45126 13072 45178
rect 13124 45126 13136 45178
rect 13188 45126 13200 45178
rect 13252 45126 14812 45178
rect 1104 45104 14812 45126
rect 1104 44634 14971 44656
rect 1104 44582 4376 44634
rect 4428 44582 4440 44634
rect 4492 44582 4504 44634
rect 4556 44582 4568 44634
rect 4620 44582 4632 44634
rect 4684 44582 7803 44634
rect 7855 44582 7867 44634
rect 7919 44582 7931 44634
rect 7983 44582 7995 44634
rect 8047 44582 8059 44634
rect 8111 44582 11230 44634
rect 11282 44582 11294 44634
rect 11346 44582 11358 44634
rect 11410 44582 11422 44634
rect 11474 44582 11486 44634
rect 11538 44582 14657 44634
rect 14709 44582 14721 44634
rect 14773 44582 14785 44634
rect 14837 44582 14849 44634
rect 14901 44582 14913 44634
rect 14965 44582 14971 44634
rect 1104 44560 14971 44582
rect 1104 44090 14812 44112
rect 1104 44038 2663 44090
rect 2715 44038 2727 44090
rect 2779 44038 2791 44090
rect 2843 44038 2855 44090
rect 2907 44038 2919 44090
rect 2971 44038 6090 44090
rect 6142 44038 6154 44090
rect 6206 44038 6218 44090
rect 6270 44038 6282 44090
rect 6334 44038 6346 44090
rect 6398 44038 9517 44090
rect 9569 44038 9581 44090
rect 9633 44038 9645 44090
rect 9697 44038 9709 44090
rect 9761 44038 9773 44090
rect 9825 44038 12944 44090
rect 12996 44038 13008 44090
rect 13060 44038 13072 44090
rect 13124 44038 13136 44090
rect 13188 44038 13200 44090
rect 13252 44038 14812 44090
rect 1104 44016 14812 44038
rect 14458 43664 14464 43716
rect 14516 43664 14522 43716
rect 1104 43546 14971 43568
rect 1104 43494 4376 43546
rect 4428 43494 4440 43546
rect 4492 43494 4504 43546
rect 4556 43494 4568 43546
rect 4620 43494 4632 43546
rect 4684 43494 7803 43546
rect 7855 43494 7867 43546
rect 7919 43494 7931 43546
rect 7983 43494 7995 43546
rect 8047 43494 8059 43546
rect 8111 43494 11230 43546
rect 11282 43494 11294 43546
rect 11346 43494 11358 43546
rect 11410 43494 11422 43546
rect 11474 43494 11486 43546
rect 11538 43494 14657 43546
rect 14709 43494 14721 43546
rect 14773 43494 14785 43546
rect 14837 43494 14849 43546
rect 14901 43494 14913 43546
rect 14965 43494 14971 43546
rect 1104 43472 14971 43494
rect 1104 43002 14812 43024
rect 1104 42950 2663 43002
rect 2715 42950 2727 43002
rect 2779 42950 2791 43002
rect 2843 42950 2855 43002
rect 2907 42950 2919 43002
rect 2971 42950 6090 43002
rect 6142 42950 6154 43002
rect 6206 42950 6218 43002
rect 6270 42950 6282 43002
rect 6334 42950 6346 43002
rect 6398 42950 9517 43002
rect 9569 42950 9581 43002
rect 9633 42950 9645 43002
rect 9697 42950 9709 43002
rect 9761 42950 9773 43002
rect 9825 42950 12944 43002
rect 12996 42950 13008 43002
rect 13060 42950 13072 43002
rect 13124 42950 13136 43002
rect 13188 42950 13200 43002
rect 13252 42950 14812 43002
rect 1104 42928 14812 42950
rect 1104 42458 14971 42480
rect 1104 42406 4376 42458
rect 4428 42406 4440 42458
rect 4492 42406 4504 42458
rect 4556 42406 4568 42458
rect 4620 42406 4632 42458
rect 4684 42406 7803 42458
rect 7855 42406 7867 42458
rect 7919 42406 7931 42458
rect 7983 42406 7995 42458
rect 8047 42406 8059 42458
rect 8111 42406 11230 42458
rect 11282 42406 11294 42458
rect 11346 42406 11358 42458
rect 11410 42406 11422 42458
rect 11474 42406 11486 42458
rect 11538 42406 14657 42458
rect 14709 42406 14721 42458
rect 14773 42406 14785 42458
rect 14837 42406 14849 42458
rect 14901 42406 14913 42458
rect 14965 42406 14971 42458
rect 1104 42384 14971 42406
rect 1104 41914 14812 41936
rect 1104 41862 2663 41914
rect 2715 41862 2727 41914
rect 2779 41862 2791 41914
rect 2843 41862 2855 41914
rect 2907 41862 2919 41914
rect 2971 41862 6090 41914
rect 6142 41862 6154 41914
rect 6206 41862 6218 41914
rect 6270 41862 6282 41914
rect 6334 41862 6346 41914
rect 6398 41862 9517 41914
rect 9569 41862 9581 41914
rect 9633 41862 9645 41914
rect 9697 41862 9709 41914
rect 9761 41862 9773 41914
rect 9825 41862 12944 41914
rect 12996 41862 13008 41914
rect 13060 41862 13072 41914
rect 13124 41862 13136 41914
rect 13188 41862 13200 41914
rect 13252 41862 14812 41914
rect 1104 41840 14812 41862
rect 1104 41370 14971 41392
rect 1104 41318 4376 41370
rect 4428 41318 4440 41370
rect 4492 41318 4504 41370
rect 4556 41318 4568 41370
rect 4620 41318 4632 41370
rect 4684 41318 7803 41370
rect 7855 41318 7867 41370
rect 7919 41318 7931 41370
rect 7983 41318 7995 41370
rect 8047 41318 8059 41370
rect 8111 41318 11230 41370
rect 11282 41318 11294 41370
rect 11346 41318 11358 41370
rect 11410 41318 11422 41370
rect 11474 41318 11486 41370
rect 11538 41318 14657 41370
rect 14709 41318 14721 41370
rect 14773 41318 14785 41370
rect 14837 41318 14849 41370
rect 14901 41318 14913 41370
rect 14965 41318 14971 41370
rect 1104 41296 14971 41318
rect 1104 40826 14812 40848
rect 1104 40774 2663 40826
rect 2715 40774 2727 40826
rect 2779 40774 2791 40826
rect 2843 40774 2855 40826
rect 2907 40774 2919 40826
rect 2971 40774 6090 40826
rect 6142 40774 6154 40826
rect 6206 40774 6218 40826
rect 6270 40774 6282 40826
rect 6334 40774 6346 40826
rect 6398 40774 9517 40826
rect 9569 40774 9581 40826
rect 9633 40774 9645 40826
rect 9697 40774 9709 40826
rect 9761 40774 9773 40826
rect 9825 40774 12944 40826
rect 12996 40774 13008 40826
rect 13060 40774 13072 40826
rect 13124 40774 13136 40826
rect 13188 40774 13200 40826
rect 13252 40774 14812 40826
rect 1104 40752 14812 40774
rect 1104 40282 14971 40304
rect 1104 40230 4376 40282
rect 4428 40230 4440 40282
rect 4492 40230 4504 40282
rect 4556 40230 4568 40282
rect 4620 40230 4632 40282
rect 4684 40230 7803 40282
rect 7855 40230 7867 40282
rect 7919 40230 7931 40282
rect 7983 40230 7995 40282
rect 8047 40230 8059 40282
rect 8111 40230 11230 40282
rect 11282 40230 11294 40282
rect 11346 40230 11358 40282
rect 11410 40230 11422 40282
rect 11474 40230 11486 40282
rect 11538 40230 14657 40282
rect 14709 40230 14721 40282
rect 14773 40230 14785 40282
rect 14837 40230 14849 40282
rect 14901 40230 14913 40282
rect 14965 40230 14971 40282
rect 1104 40208 14971 40230
rect 1104 39738 14812 39760
rect 1104 39686 2663 39738
rect 2715 39686 2727 39738
rect 2779 39686 2791 39738
rect 2843 39686 2855 39738
rect 2907 39686 2919 39738
rect 2971 39686 6090 39738
rect 6142 39686 6154 39738
rect 6206 39686 6218 39738
rect 6270 39686 6282 39738
rect 6334 39686 6346 39738
rect 6398 39686 9517 39738
rect 9569 39686 9581 39738
rect 9633 39686 9645 39738
rect 9697 39686 9709 39738
rect 9761 39686 9773 39738
rect 9825 39686 12944 39738
rect 12996 39686 13008 39738
rect 13060 39686 13072 39738
rect 13124 39686 13136 39738
rect 13188 39686 13200 39738
rect 13252 39686 14812 39738
rect 1104 39664 14812 39686
rect 1104 39194 14971 39216
rect 1104 39142 4376 39194
rect 4428 39142 4440 39194
rect 4492 39142 4504 39194
rect 4556 39142 4568 39194
rect 4620 39142 4632 39194
rect 4684 39142 7803 39194
rect 7855 39142 7867 39194
rect 7919 39142 7931 39194
rect 7983 39142 7995 39194
rect 8047 39142 8059 39194
rect 8111 39142 11230 39194
rect 11282 39142 11294 39194
rect 11346 39142 11358 39194
rect 11410 39142 11422 39194
rect 11474 39142 11486 39194
rect 11538 39142 14657 39194
rect 14709 39142 14721 39194
rect 14773 39142 14785 39194
rect 14837 39142 14849 39194
rect 14901 39142 14913 39194
rect 14965 39142 14971 39194
rect 1104 39120 14971 39142
rect 1104 38650 14812 38672
rect 1104 38598 2663 38650
rect 2715 38598 2727 38650
rect 2779 38598 2791 38650
rect 2843 38598 2855 38650
rect 2907 38598 2919 38650
rect 2971 38598 6090 38650
rect 6142 38598 6154 38650
rect 6206 38598 6218 38650
rect 6270 38598 6282 38650
rect 6334 38598 6346 38650
rect 6398 38598 9517 38650
rect 9569 38598 9581 38650
rect 9633 38598 9645 38650
rect 9697 38598 9709 38650
rect 9761 38598 9773 38650
rect 9825 38598 12944 38650
rect 12996 38598 13008 38650
rect 13060 38598 13072 38650
rect 13124 38598 13136 38650
rect 13188 38598 13200 38650
rect 13252 38598 14812 38650
rect 1104 38576 14812 38598
rect 1104 38106 14971 38128
rect 1104 38054 4376 38106
rect 4428 38054 4440 38106
rect 4492 38054 4504 38106
rect 4556 38054 4568 38106
rect 4620 38054 4632 38106
rect 4684 38054 7803 38106
rect 7855 38054 7867 38106
rect 7919 38054 7931 38106
rect 7983 38054 7995 38106
rect 8047 38054 8059 38106
rect 8111 38054 11230 38106
rect 11282 38054 11294 38106
rect 11346 38054 11358 38106
rect 11410 38054 11422 38106
rect 11474 38054 11486 38106
rect 11538 38054 14657 38106
rect 14709 38054 14721 38106
rect 14773 38054 14785 38106
rect 14837 38054 14849 38106
rect 14901 38054 14913 38106
rect 14965 38054 14971 38106
rect 1104 38032 14971 38054
rect 1104 37562 14812 37584
rect 1104 37510 2663 37562
rect 2715 37510 2727 37562
rect 2779 37510 2791 37562
rect 2843 37510 2855 37562
rect 2907 37510 2919 37562
rect 2971 37510 6090 37562
rect 6142 37510 6154 37562
rect 6206 37510 6218 37562
rect 6270 37510 6282 37562
rect 6334 37510 6346 37562
rect 6398 37510 9517 37562
rect 9569 37510 9581 37562
rect 9633 37510 9645 37562
rect 9697 37510 9709 37562
rect 9761 37510 9773 37562
rect 9825 37510 12944 37562
rect 12996 37510 13008 37562
rect 13060 37510 13072 37562
rect 13124 37510 13136 37562
rect 13188 37510 13200 37562
rect 13252 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14971 37040
rect 1104 36966 4376 37018
rect 4428 36966 4440 37018
rect 4492 36966 4504 37018
rect 4556 36966 4568 37018
rect 4620 36966 4632 37018
rect 4684 36966 7803 37018
rect 7855 36966 7867 37018
rect 7919 36966 7931 37018
rect 7983 36966 7995 37018
rect 8047 36966 8059 37018
rect 8111 36966 11230 37018
rect 11282 36966 11294 37018
rect 11346 36966 11358 37018
rect 11410 36966 11422 37018
rect 11474 36966 11486 37018
rect 11538 36966 14657 37018
rect 14709 36966 14721 37018
rect 14773 36966 14785 37018
rect 14837 36966 14849 37018
rect 14901 36966 14913 37018
rect 14965 36966 14971 37018
rect 1104 36944 14971 36966
rect 1104 36474 14812 36496
rect 1104 36422 2663 36474
rect 2715 36422 2727 36474
rect 2779 36422 2791 36474
rect 2843 36422 2855 36474
rect 2907 36422 2919 36474
rect 2971 36422 6090 36474
rect 6142 36422 6154 36474
rect 6206 36422 6218 36474
rect 6270 36422 6282 36474
rect 6334 36422 6346 36474
rect 6398 36422 9517 36474
rect 9569 36422 9581 36474
rect 9633 36422 9645 36474
rect 9697 36422 9709 36474
rect 9761 36422 9773 36474
rect 9825 36422 12944 36474
rect 12996 36422 13008 36474
rect 13060 36422 13072 36474
rect 13124 36422 13136 36474
rect 13188 36422 13200 36474
rect 13252 36422 14812 36474
rect 1104 36400 14812 36422
rect 14458 35980 14464 36032
rect 14516 35980 14522 36032
rect 1104 35930 14971 35952
rect 1104 35878 4376 35930
rect 4428 35878 4440 35930
rect 4492 35878 4504 35930
rect 4556 35878 4568 35930
rect 4620 35878 4632 35930
rect 4684 35878 7803 35930
rect 7855 35878 7867 35930
rect 7919 35878 7931 35930
rect 7983 35878 7995 35930
rect 8047 35878 8059 35930
rect 8111 35878 11230 35930
rect 11282 35878 11294 35930
rect 11346 35878 11358 35930
rect 11410 35878 11422 35930
rect 11474 35878 11486 35930
rect 11538 35878 14657 35930
rect 14709 35878 14721 35930
rect 14773 35878 14785 35930
rect 14837 35878 14849 35930
rect 14901 35878 14913 35930
rect 14965 35878 14971 35930
rect 1104 35856 14971 35878
rect 1104 35386 14812 35408
rect 1104 35334 2663 35386
rect 2715 35334 2727 35386
rect 2779 35334 2791 35386
rect 2843 35334 2855 35386
rect 2907 35334 2919 35386
rect 2971 35334 6090 35386
rect 6142 35334 6154 35386
rect 6206 35334 6218 35386
rect 6270 35334 6282 35386
rect 6334 35334 6346 35386
rect 6398 35334 9517 35386
rect 9569 35334 9581 35386
rect 9633 35334 9645 35386
rect 9697 35334 9709 35386
rect 9761 35334 9773 35386
rect 9825 35334 12944 35386
rect 12996 35334 13008 35386
rect 13060 35334 13072 35386
rect 13124 35334 13136 35386
rect 13188 35334 13200 35386
rect 13252 35334 14812 35386
rect 1104 35312 14812 35334
rect 1104 34842 14971 34864
rect 1104 34790 4376 34842
rect 4428 34790 4440 34842
rect 4492 34790 4504 34842
rect 4556 34790 4568 34842
rect 4620 34790 4632 34842
rect 4684 34790 7803 34842
rect 7855 34790 7867 34842
rect 7919 34790 7931 34842
rect 7983 34790 7995 34842
rect 8047 34790 8059 34842
rect 8111 34790 11230 34842
rect 11282 34790 11294 34842
rect 11346 34790 11358 34842
rect 11410 34790 11422 34842
rect 11474 34790 11486 34842
rect 11538 34790 14657 34842
rect 14709 34790 14721 34842
rect 14773 34790 14785 34842
rect 14837 34790 14849 34842
rect 14901 34790 14913 34842
rect 14965 34790 14971 34842
rect 1104 34768 14971 34790
rect 1104 34298 14812 34320
rect 1104 34246 2663 34298
rect 2715 34246 2727 34298
rect 2779 34246 2791 34298
rect 2843 34246 2855 34298
rect 2907 34246 2919 34298
rect 2971 34246 6090 34298
rect 6142 34246 6154 34298
rect 6206 34246 6218 34298
rect 6270 34246 6282 34298
rect 6334 34246 6346 34298
rect 6398 34246 9517 34298
rect 9569 34246 9581 34298
rect 9633 34246 9645 34298
rect 9697 34246 9709 34298
rect 9761 34246 9773 34298
rect 9825 34246 12944 34298
rect 12996 34246 13008 34298
rect 13060 34246 13072 34298
rect 13124 34246 13136 34298
rect 13188 34246 13200 34298
rect 13252 34246 14812 34298
rect 1104 34224 14812 34246
rect 1104 33754 14971 33776
rect 1104 33702 4376 33754
rect 4428 33702 4440 33754
rect 4492 33702 4504 33754
rect 4556 33702 4568 33754
rect 4620 33702 4632 33754
rect 4684 33702 7803 33754
rect 7855 33702 7867 33754
rect 7919 33702 7931 33754
rect 7983 33702 7995 33754
rect 8047 33702 8059 33754
rect 8111 33702 11230 33754
rect 11282 33702 11294 33754
rect 11346 33702 11358 33754
rect 11410 33702 11422 33754
rect 11474 33702 11486 33754
rect 11538 33702 14657 33754
rect 14709 33702 14721 33754
rect 14773 33702 14785 33754
rect 14837 33702 14849 33754
rect 14901 33702 14913 33754
rect 14965 33702 14971 33754
rect 1104 33680 14971 33702
rect 1104 33210 14812 33232
rect 1104 33158 2663 33210
rect 2715 33158 2727 33210
rect 2779 33158 2791 33210
rect 2843 33158 2855 33210
rect 2907 33158 2919 33210
rect 2971 33158 6090 33210
rect 6142 33158 6154 33210
rect 6206 33158 6218 33210
rect 6270 33158 6282 33210
rect 6334 33158 6346 33210
rect 6398 33158 9517 33210
rect 9569 33158 9581 33210
rect 9633 33158 9645 33210
rect 9697 33158 9709 33210
rect 9761 33158 9773 33210
rect 9825 33158 12944 33210
rect 12996 33158 13008 33210
rect 13060 33158 13072 33210
rect 13124 33158 13136 33210
rect 13188 33158 13200 33210
rect 13252 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14971 32688
rect 1104 32614 4376 32666
rect 4428 32614 4440 32666
rect 4492 32614 4504 32666
rect 4556 32614 4568 32666
rect 4620 32614 4632 32666
rect 4684 32614 7803 32666
rect 7855 32614 7867 32666
rect 7919 32614 7931 32666
rect 7983 32614 7995 32666
rect 8047 32614 8059 32666
rect 8111 32614 11230 32666
rect 11282 32614 11294 32666
rect 11346 32614 11358 32666
rect 11410 32614 11422 32666
rect 11474 32614 11486 32666
rect 11538 32614 14657 32666
rect 14709 32614 14721 32666
rect 14773 32614 14785 32666
rect 14837 32614 14849 32666
rect 14901 32614 14913 32666
rect 14965 32614 14971 32666
rect 1104 32592 14971 32614
rect 1104 32122 14812 32144
rect 1104 32070 2663 32122
rect 2715 32070 2727 32122
rect 2779 32070 2791 32122
rect 2843 32070 2855 32122
rect 2907 32070 2919 32122
rect 2971 32070 6090 32122
rect 6142 32070 6154 32122
rect 6206 32070 6218 32122
rect 6270 32070 6282 32122
rect 6334 32070 6346 32122
rect 6398 32070 9517 32122
rect 9569 32070 9581 32122
rect 9633 32070 9645 32122
rect 9697 32070 9709 32122
rect 9761 32070 9773 32122
rect 9825 32070 12944 32122
rect 12996 32070 13008 32122
rect 13060 32070 13072 32122
rect 13124 32070 13136 32122
rect 13188 32070 13200 32122
rect 13252 32070 14812 32122
rect 1104 32048 14812 32070
rect 1104 31578 14971 31600
rect 1104 31526 4376 31578
rect 4428 31526 4440 31578
rect 4492 31526 4504 31578
rect 4556 31526 4568 31578
rect 4620 31526 4632 31578
rect 4684 31526 7803 31578
rect 7855 31526 7867 31578
rect 7919 31526 7931 31578
rect 7983 31526 7995 31578
rect 8047 31526 8059 31578
rect 8111 31526 11230 31578
rect 11282 31526 11294 31578
rect 11346 31526 11358 31578
rect 11410 31526 11422 31578
rect 11474 31526 11486 31578
rect 11538 31526 14657 31578
rect 14709 31526 14721 31578
rect 14773 31526 14785 31578
rect 14837 31526 14849 31578
rect 14901 31526 14913 31578
rect 14965 31526 14971 31578
rect 1104 31504 14971 31526
rect 1104 31034 14812 31056
rect 1104 30982 2663 31034
rect 2715 30982 2727 31034
rect 2779 30982 2791 31034
rect 2843 30982 2855 31034
rect 2907 30982 2919 31034
rect 2971 30982 6090 31034
rect 6142 30982 6154 31034
rect 6206 30982 6218 31034
rect 6270 30982 6282 31034
rect 6334 30982 6346 31034
rect 6398 30982 9517 31034
rect 9569 30982 9581 31034
rect 9633 30982 9645 31034
rect 9697 30982 9709 31034
rect 9761 30982 9773 31034
rect 9825 30982 12944 31034
rect 12996 30982 13008 31034
rect 13060 30982 13072 31034
rect 13124 30982 13136 31034
rect 13188 30982 13200 31034
rect 13252 30982 14812 31034
rect 1104 30960 14812 30982
rect 1104 30490 14971 30512
rect 1104 30438 4376 30490
rect 4428 30438 4440 30490
rect 4492 30438 4504 30490
rect 4556 30438 4568 30490
rect 4620 30438 4632 30490
rect 4684 30438 7803 30490
rect 7855 30438 7867 30490
rect 7919 30438 7931 30490
rect 7983 30438 7995 30490
rect 8047 30438 8059 30490
rect 8111 30438 11230 30490
rect 11282 30438 11294 30490
rect 11346 30438 11358 30490
rect 11410 30438 11422 30490
rect 11474 30438 11486 30490
rect 11538 30438 14657 30490
rect 14709 30438 14721 30490
rect 14773 30438 14785 30490
rect 14837 30438 14849 30490
rect 14901 30438 14913 30490
rect 14965 30438 14971 30490
rect 1104 30416 14971 30438
rect 1104 29946 14812 29968
rect 1104 29894 2663 29946
rect 2715 29894 2727 29946
rect 2779 29894 2791 29946
rect 2843 29894 2855 29946
rect 2907 29894 2919 29946
rect 2971 29894 6090 29946
rect 6142 29894 6154 29946
rect 6206 29894 6218 29946
rect 6270 29894 6282 29946
rect 6334 29894 6346 29946
rect 6398 29894 9517 29946
rect 9569 29894 9581 29946
rect 9633 29894 9645 29946
rect 9697 29894 9709 29946
rect 9761 29894 9773 29946
rect 9825 29894 12944 29946
rect 12996 29894 13008 29946
rect 13060 29894 13072 29946
rect 13124 29894 13136 29946
rect 13188 29894 13200 29946
rect 13252 29894 14812 29946
rect 1104 29872 14812 29894
rect 1104 29402 14971 29424
rect 1104 29350 4376 29402
rect 4428 29350 4440 29402
rect 4492 29350 4504 29402
rect 4556 29350 4568 29402
rect 4620 29350 4632 29402
rect 4684 29350 7803 29402
rect 7855 29350 7867 29402
rect 7919 29350 7931 29402
rect 7983 29350 7995 29402
rect 8047 29350 8059 29402
rect 8111 29350 11230 29402
rect 11282 29350 11294 29402
rect 11346 29350 11358 29402
rect 11410 29350 11422 29402
rect 11474 29350 11486 29402
rect 11538 29350 14657 29402
rect 14709 29350 14721 29402
rect 14773 29350 14785 29402
rect 14837 29350 14849 29402
rect 14901 29350 14913 29402
rect 14965 29350 14971 29402
rect 1104 29328 14971 29350
rect 1104 28858 14812 28880
rect 1104 28806 2663 28858
rect 2715 28806 2727 28858
rect 2779 28806 2791 28858
rect 2843 28806 2855 28858
rect 2907 28806 2919 28858
rect 2971 28806 6090 28858
rect 6142 28806 6154 28858
rect 6206 28806 6218 28858
rect 6270 28806 6282 28858
rect 6334 28806 6346 28858
rect 6398 28806 9517 28858
rect 9569 28806 9581 28858
rect 9633 28806 9645 28858
rect 9697 28806 9709 28858
rect 9761 28806 9773 28858
rect 9825 28806 12944 28858
rect 12996 28806 13008 28858
rect 13060 28806 13072 28858
rect 13124 28806 13136 28858
rect 13188 28806 13200 28858
rect 13252 28806 14812 28858
rect 1104 28784 14812 28806
rect 1104 28314 14971 28336
rect 1104 28262 4376 28314
rect 4428 28262 4440 28314
rect 4492 28262 4504 28314
rect 4556 28262 4568 28314
rect 4620 28262 4632 28314
rect 4684 28262 7803 28314
rect 7855 28262 7867 28314
rect 7919 28262 7931 28314
rect 7983 28262 7995 28314
rect 8047 28262 8059 28314
rect 8111 28262 11230 28314
rect 11282 28262 11294 28314
rect 11346 28262 11358 28314
rect 11410 28262 11422 28314
rect 11474 28262 11486 28314
rect 11538 28262 14657 28314
rect 14709 28262 14721 28314
rect 14773 28262 14785 28314
rect 14837 28262 14849 28314
rect 14901 28262 14913 28314
rect 14965 28262 14971 28314
rect 1104 28240 14971 28262
rect 14458 27956 14464 28008
rect 14516 27956 14522 28008
rect 1104 27770 14812 27792
rect 1104 27718 2663 27770
rect 2715 27718 2727 27770
rect 2779 27718 2791 27770
rect 2843 27718 2855 27770
rect 2907 27718 2919 27770
rect 2971 27718 6090 27770
rect 6142 27718 6154 27770
rect 6206 27718 6218 27770
rect 6270 27718 6282 27770
rect 6334 27718 6346 27770
rect 6398 27718 9517 27770
rect 9569 27718 9581 27770
rect 9633 27718 9645 27770
rect 9697 27718 9709 27770
rect 9761 27718 9773 27770
rect 9825 27718 12944 27770
rect 12996 27718 13008 27770
rect 13060 27718 13072 27770
rect 13124 27718 13136 27770
rect 13188 27718 13200 27770
rect 13252 27718 14812 27770
rect 1104 27696 14812 27718
rect 1104 27226 14971 27248
rect 1104 27174 4376 27226
rect 4428 27174 4440 27226
rect 4492 27174 4504 27226
rect 4556 27174 4568 27226
rect 4620 27174 4632 27226
rect 4684 27174 7803 27226
rect 7855 27174 7867 27226
rect 7919 27174 7931 27226
rect 7983 27174 7995 27226
rect 8047 27174 8059 27226
rect 8111 27174 11230 27226
rect 11282 27174 11294 27226
rect 11346 27174 11358 27226
rect 11410 27174 11422 27226
rect 11474 27174 11486 27226
rect 11538 27174 14657 27226
rect 14709 27174 14721 27226
rect 14773 27174 14785 27226
rect 14837 27174 14849 27226
rect 14901 27174 14913 27226
rect 14965 27174 14971 27226
rect 1104 27152 14971 27174
rect 1104 26682 14812 26704
rect 1104 26630 2663 26682
rect 2715 26630 2727 26682
rect 2779 26630 2791 26682
rect 2843 26630 2855 26682
rect 2907 26630 2919 26682
rect 2971 26630 6090 26682
rect 6142 26630 6154 26682
rect 6206 26630 6218 26682
rect 6270 26630 6282 26682
rect 6334 26630 6346 26682
rect 6398 26630 9517 26682
rect 9569 26630 9581 26682
rect 9633 26630 9645 26682
rect 9697 26630 9709 26682
rect 9761 26630 9773 26682
rect 9825 26630 12944 26682
rect 12996 26630 13008 26682
rect 13060 26630 13072 26682
rect 13124 26630 13136 26682
rect 13188 26630 13200 26682
rect 13252 26630 14812 26682
rect 1104 26608 14812 26630
rect 1104 26138 14971 26160
rect 1104 26086 4376 26138
rect 4428 26086 4440 26138
rect 4492 26086 4504 26138
rect 4556 26086 4568 26138
rect 4620 26086 4632 26138
rect 4684 26086 7803 26138
rect 7855 26086 7867 26138
rect 7919 26086 7931 26138
rect 7983 26086 7995 26138
rect 8047 26086 8059 26138
rect 8111 26086 11230 26138
rect 11282 26086 11294 26138
rect 11346 26086 11358 26138
rect 11410 26086 11422 26138
rect 11474 26086 11486 26138
rect 11538 26086 14657 26138
rect 14709 26086 14721 26138
rect 14773 26086 14785 26138
rect 14837 26086 14849 26138
rect 14901 26086 14913 26138
rect 14965 26086 14971 26138
rect 1104 26064 14971 26086
rect 1104 25594 14812 25616
rect 1104 25542 2663 25594
rect 2715 25542 2727 25594
rect 2779 25542 2791 25594
rect 2843 25542 2855 25594
rect 2907 25542 2919 25594
rect 2971 25542 6090 25594
rect 6142 25542 6154 25594
rect 6206 25542 6218 25594
rect 6270 25542 6282 25594
rect 6334 25542 6346 25594
rect 6398 25542 9517 25594
rect 9569 25542 9581 25594
rect 9633 25542 9645 25594
rect 9697 25542 9709 25594
rect 9761 25542 9773 25594
rect 9825 25542 12944 25594
rect 12996 25542 13008 25594
rect 13060 25542 13072 25594
rect 13124 25542 13136 25594
rect 13188 25542 13200 25594
rect 13252 25542 14812 25594
rect 1104 25520 14812 25542
rect 1104 25050 14971 25072
rect 1104 24998 4376 25050
rect 4428 24998 4440 25050
rect 4492 24998 4504 25050
rect 4556 24998 4568 25050
rect 4620 24998 4632 25050
rect 4684 24998 7803 25050
rect 7855 24998 7867 25050
rect 7919 24998 7931 25050
rect 7983 24998 7995 25050
rect 8047 24998 8059 25050
rect 8111 24998 11230 25050
rect 11282 24998 11294 25050
rect 11346 24998 11358 25050
rect 11410 24998 11422 25050
rect 11474 24998 11486 25050
rect 11538 24998 14657 25050
rect 14709 24998 14721 25050
rect 14773 24998 14785 25050
rect 14837 24998 14849 25050
rect 14901 24998 14913 25050
rect 14965 24998 14971 25050
rect 1104 24976 14971 24998
rect 1104 24506 14812 24528
rect 1104 24454 2663 24506
rect 2715 24454 2727 24506
rect 2779 24454 2791 24506
rect 2843 24454 2855 24506
rect 2907 24454 2919 24506
rect 2971 24454 6090 24506
rect 6142 24454 6154 24506
rect 6206 24454 6218 24506
rect 6270 24454 6282 24506
rect 6334 24454 6346 24506
rect 6398 24454 9517 24506
rect 9569 24454 9581 24506
rect 9633 24454 9645 24506
rect 9697 24454 9709 24506
rect 9761 24454 9773 24506
rect 9825 24454 12944 24506
rect 12996 24454 13008 24506
rect 13060 24454 13072 24506
rect 13124 24454 13136 24506
rect 13188 24454 13200 24506
rect 13252 24454 14812 24506
rect 1104 24432 14812 24454
rect 1104 23962 14971 23984
rect 1104 23910 4376 23962
rect 4428 23910 4440 23962
rect 4492 23910 4504 23962
rect 4556 23910 4568 23962
rect 4620 23910 4632 23962
rect 4684 23910 7803 23962
rect 7855 23910 7867 23962
rect 7919 23910 7931 23962
rect 7983 23910 7995 23962
rect 8047 23910 8059 23962
rect 8111 23910 11230 23962
rect 11282 23910 11294 23962
rect 11346 23910 11358 23962
rect 11410 23910 11422 23962
rect 11474 23910 11486 23962
rect 11538 23910 14657 23962
rect 14709 23910 14721 23962
rect 14773 23910 14785 23962
rect 14837 23910 14849 23962
rect 14901 23910 14913 23962
rect 14965 23910 14971 23962
rect 1104 23888 14971 23910
rect 1104 23418 14812 23440
rect 1104 23366 2663 23418
rect 2715 23366 2727 23418
rect 2779 23366 2791 23418
rect 2843 23366 2855 23418
rect 2907 23366 2919 23418
rect 2971 23366 6090 23418
rect 6142 23366 6154 23418
rect 6206 23366 6218 23418
rect 6270 23366 6282 23418
rect 6334 23366 6346 23418
rect 6398 23366 9517 23418
rect 9569 23366 9581 23418
rect 9633 23366 9645 23418
rect 9697 23366 9709 23418
rect 9761 23366 9773 23418
rect 9825 23366 12944 23418
rect 12996 23366 13008 23418
rect 13060 23366 13072 23418
rect 13124 23366 13136 23418
rect 13188 23366 13200 23418
rect 13252 23366 14812 23418
rect 1104 23344 14812 23366
rect 1104 22874 14971 22896
rect 1104 22822 4376 22874
rect 4428 22822 4440 22874
rect 4492 22822 4504 22874
rect 4556 22822 4568 22874
rect 4620 22822 4632 22874
rect 4684 22822 7803 22874
rect 7855 22822 7867 22874
rect 7919 22822 7931 22874
rect 7983 22822 7995 22874
rect 8047 22822 8059 22874
rect 8111 22822 11230 22874
rect 11282 22822 11294 22874
rect 11346 22822 11358 22874
rect 11410 22822 11422 22874
rect 11474 22822 11486 22874
rect 11538 22822 14657 22874
rect 14709 22822 14721 22874
rect 14773 22822 14785 22874
rect 14837 22822 14849 22874
rect 14901 22822 14913 22874
rect 14965 22822 14971 22874
rect 1104 22800 14971 22822
rect 1104 22330 14812 22352
rect 1104 22278 2663 22330
rect 2715 22278 2727 22330
rect 2779 22278 2791 22330
rect 2843 22278 2855 22330
rect 2907 22278 2919 22330
rect 2971 22278 6090 22330
rect 6142 22278 6154 22330
rect 6206 22278 6218 22330
rect 6270 22278 6282 22330
rect 6334 22278 6346 22330
rect 6398 22278 9517 22330
rect 9569 22278 9581 22330
rect 9633 22278 9645 22330
rect 9697 22278 9709 22330
rect 9761 22278 9773 22330
rect 9825 22278 12944 22330
rect 12996 22278 13008 22330
rect 13060 22278 13072 22330
rect 13124 22278 13136 22330
rect 13188 22278 13200 22330
rect 13252 22278 14812 22330
rect 1104 22256 14812 22278
rect 1104 21786 14971 21808
rect 1104 21734 4376 21786
rect 4428 21734 4440 21786
rect 4492 21734 4504 21786
rect 4556 21734 4568 21786
rect 4620 21734 4632 21786
rect 4684 21734 7803 21786
rect 7855 21734 7867 21786
rect 7919 21734 7931 21786
rect 7983 21734 7995 21786
rect 8047 21734 8059 21786
rect 8111 21734 11230 21786
rect 11282 21734 11294 21786
rect 11346 21734 11358 21786
rect 11410 21734 11422 21786
rect 11474 21734 11486 21786
rect 11538 21734 14657 21786
rect 14709 21734 14721 21786
rect 14773 21734 14785 21786
rect 14837 21734 14849 21786
rect 14901 21734 14913 21786
rect 14965 21734 14971 21786
rect 1104 21712 14971 21734
rect 1104 21242 14812 21264
rect 1104 21190 2663 21242
rect 2715 21190 2727 21242
rect 2779 21190 2791 21242
rect 2843 21190 2855 21242
rect 2907 21190 2919 21242
rect 2971 21190 6090 21242
rect 6142 21190 6154 21242
rect 6206 21190 6218 21242
rect 6270 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 9517 21242
rect 9569 21190 9581 21242
rect 9633 21190 9645 21242
rect 9697 21190 9709 21242
rect 9761 21190 9773 21242
rect 9825 21190 12944 21242
rect 12996 21190 13008 21242
rect 13060 21190 13072 21242
rect 13124 21190 13136 21242
rect 13188 21190 13200 21242
rect 13252 21190 14812 21242
rect 1104 21168 14812 21190
rect 1104 20698 14971 20720
rect 1104 20646 4376 20698
rect 4428 20646 4440 20698
rect 4492 20646 4504 20698
rect 4556 20646 4568 20698
rect 4620 20646 4632 20698
rect 4684 20646 7803 20698
rect 7855 20646 7867 20698
rect 7919 20646 7931 20698
rect 7983 20646 7995 20698
rect 8047 20646 8059 20698
rect 8111 20646 11230 20698
rect 11282 20646 11294 20698
rect 11346 20646 11358 20698
rect 11410 20646 11422 20698
rect 11474 20646 11486 20698
rect 11538 20646 14657 20698
rect 14709 20646 14721 20698
rect 14773 20646 14785 20698
rect 14837 20646 14849 20698
rect 14901 20646 14913 20698
rect 14965 20646 14971 20698
rect 1104 20624 14971 20646
rect 14458 20340 14464 20392
rect 14516 20340 14522 20392
rect 1104 20154 14812 20176
rect 1104 20102 2663 20154
rect 2715 20102 2727 20154
rect 2779 20102 2791 20154
rect 2843 20102 2855 20154
rect 2907 20102 2919 20154
rect 2971 20102 6090 20154
rect 6142 20102 6154 20154
rect 6206 20102 6218 20154
rect 6270 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 9517 20154
rect 9569 20102 9581 20154
rect 9633 20102 9645 20154
rect 9697 20102 9709 20154
rect 9761 20102 9773 20154
rect 9825 20102 12944 20154
rect 12996 20102 13008 20154
rect 13060 20102 13072 20154
rect 13124 20102 13136 20154
rect 13188 20102 13200 20154
rect 13252 20102 14812 20154
rect 1104 20080 14812 20102
rect 1104 19610 14971 19632
rect 1104 19558 4376 19610
rect 4428 19558 4440 19610
rect 4492 19558 4504 19610
rect 4556 19558 4568 19610
rect 4620 19558 4632 19610
rect 4684 19558 7803 19610
rect 7855 19558 7867 19610
rect 7919 19558 7931 19610
rect 7983 19558 7995 19610
rect 8047 19558 8059 19610
rect 8111 19558 11230 19610
rect 11282 19558 11294 19610
rect 11346 19558 11358 19610
rect 11410 19558 11422 19610
rect 11474 19558 11486 19610
rect 11538 19558 14657 19610
rect 14709 19558 14721 19610
rect 14773 19558 14785 19610
rect 14837 19558 14849 19610
rect 14901 19558 14913 19610
rect 14965 19558 14971 19610
rect 1104 19536 14971 19558
rect 1104 19066 14812 19088
rect 1104 19014 2663 19066
rect 2715 19014 2727 19066
rect 2779 19014 2791 19066
rect 2843 19014 2855 19066
rect 2907 19014 2919 19066
rect 2971 19014 6090 19066
rect 6142 19014 6154 19066
rect 6206 19014 6218 19066
rect 6270 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 9517 19066
rect 9569 19014 9581 19066
rect 9633 19014 9645 19066
rect 9697 19014 9709 19066
rect 9761 19014 9773 19066
rect 9825 19014 12944 19066
rect 12996 19014 13008 19066
rect 13060 19014 13072 19066
rect 13124 19014 13136 19066
rect 13188 19014 13200 19066
rect 13252 19014 14812 19066
rect 1104 18992 14812 19014
rect 1104 18522 14971 18544
rect 1104 18470 4376 18522
rect 4428 18470 4440 18522
rect 4492 18470 4504 18522
rect 4556 18470 4568 18522
rect 4620 18470 4632 18522
rect 4684 18470 7803 18522
rect 7855 18470 7867 18522
rect 7919 18470 7931 18522
rect 7983 18470 7995 18522
rect 8047 18470 8059 18522
rect 8111 18470 11230 18522
rect 11282 18470 11294 18522
rect 11346 18470 11358 18522
rect 11410 18470 11422 18522
rect 11474 18470 11486 18522
rect 11538 18470 14657 18522
rect 14709 18470 14721 18522
rect 14773 18470 14785 18522
rect 14837 18470 14849 18522
rect 14901 18470 14913 18522
rect 14965 18470 14971 18522
rect 1104 18448 14971 18470
rect 1104 17978 14812 18000
rect 1104 17926 2663 17978
rect 2715 17926 2727 17978
rect 2779 17926 2791 17978
rect 2843 17926 2855 17978
rect 2907 17926 2919 17978
rect 2971 17926 6090 17978
rect 6142 17926 6154 17978
rect 6206 17926 6218 17978
rect 6270 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 9517 17978
rect 9569 17926 9581 17978
rect 9633 17926 9645 17978
rect 9697 17926 9709 17978
rect 9761 17926 9773 17978
rect 9825 17926 12944 17978
rect 12996 17926 13008 17978
rect 13060 17926 13072 17978
rect 13124 17926 13136 17978
rect 13188 17926 13200 17978
rect 13252 17926 14812 17978
rect 1104 17904 14812 17926
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 14458 12112 14464 12164
rect 14516 12112 14522 12164
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 14458 4428 14464 4480
rect 14516 4428 14522 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
<< via1 >>
rect 4376 45670 4428 45722
rect 4440 45670 4492 45722
rect 4504 45670 4556 45722
rect 4568 45670 4620 45722
rect 4632 45670 4684 45722
rect 7803 45670 7855 45722
rect 7867 45670 7919 45722
rect 7931 45670 7983 45722
rect 7995 45670 8047 45722
rect 8059 45670 8111 45722
rect 11230 45670 11282 45722
rect 11294 45670 11346 45722
rect 11358 45670 11410 45722
rect 11422 45670 11474 45722
rect 11486 45670 11538 45722
rect 14657 45670 14709 45722
rect 14721 45670 14773 45722
rect 14785 45670 14837 45722
rect 14849 45670 14901 45722
rect 14913 45670 14965 45722
rect 2663 45126 2715 45178
rect 2727 45126 2779 45178
rect 2791 45126 2843 45178
rect 2855 45126 2907 45178
rect 2919 45126 2971 45178
rect 6090 45126 6142 45178
rect 6154 45126 6206 45178
rect 6218 45126 6270 45178
rect 6282 45126 6334 45178
rect 6346 45126 6398 45178
rect 9517 45126 9569 45178
rect 9581 45126 9633 45178
rect 9645 45126 9697 45178
rect 9709 45126 9761 45178
rect 9773 45126 9825 45178
rect 12944 45126 12996 45178
rect 13008 45126 13060 45178
rect 13072 45126 13124 45178
rect 13136 45126 13188 45178
rect 13200 45126 13252 45178
rect 4376 44582 4428 44634
rect 4440 44582 4492 44634
rect 4504 44582 4556 44634
rect 4568 44582 4620 44634
rect 4632 44582 4684 44634
rect 7803 44582 7855 44634
rect 7867 44582 7919 44634
rect 7931 44582 7983 44634
rect 7995 44582 8047 44634
rect 8059 44582 8111 44634
rect 11230 44582 11282 44634
rect 11294 44582 11346 44634
rect 11358 44582 11410 44634
rect 11422 44582 11474 44634
rect 11486 44582 11538 44634
rect 14657 44582 14709 44634
rect 14721 44582 14773 44634
rect 14785 44582 14837 44634
rect 14849 44582 14901 44634
rect 14913 44582 14965 44634
rect 2663 44038 2715 44090
rect 2727 44038 2779 44090
rect 2791 44038 2843 44090
rect 2855 44038 2907 44090
rect 2919 44038 2971 44090
rect 6090 44038 6142 44090
rect 6154 44038 6206 44090
rect 6218 44038 6270 44090
rect 6282 44038 6334 44090
rect 6346 44038 6398 44090
rect 9517 44038 9569 44090
rect 9581 44038 9633 44090
rect 9645 44038 9697 44090
rect 9709 44038 9761 44090
rect 9773 44038 9825 44090
rect 12944 44038 12996 44090
rect 13008 44038 13060 44090
rect 13072 44038 13124 44090
rect 13136 44038 13188 44090
rect 13200 44038 13252 44090
rect 14464 43707 14516 43716
rect 14464 43673 14473 43707
rect 14473 43673 14507 43707
rect 14507 43673 14516 43707
rect 14464 43664 14516 43673
rect 4376 43494 4428 43546
rect 4440 43494 4492 43546
rect 4504 43494 4556 43546
rect 4568 43494 4620 43546
rect 4632 43494 4684 43546
rect 7803 43494 7855 43546
rect 7867 43494 7919 43546
rect 7931 43494 7983 43546
rect 7995 43494 8047 43546
rect 8059 43494 8111 43546
rect 11230 43494 11282 43546
rect 11294 43494 11346 43546
rect 11358 43494 11410 43546
rect 11422 43494 11474 43546
rect 11486 43494 11538 43546
rect 14657 43494 14709 43546
rect 14721 43494 14773 43546
rect 14785 43494 14837 43546
rect 14849 43494 14901 43546
rect 14913 43494 14965 43546
rect 2663 42950 2715 43002
rect 2727 42950 2779 43002
rect 2791 42950 2843 43002
rect 2855 42950 2907 43002
rect 2919 42950 2971 43002
rect 6090 42950 6142 43002
rect 6154 42950 6206 43002
rect 6218 42950 6270 43002
rect 6282 42950 6334 43002
rect 6346 42950 6398 43002
rect 9517 42950 9569 43002
rect 9581 42950 9633 43002
rect 9645 42950 9697 43002
rect 9709 42950 9761 43002
rect 9773 42950 9825 43002
rect 12944 42950 12996 43002
rect 13008 42950 13060 43002
rect 13072 42950 13124 43002
rect 13136 42950 13188 43002
rect 13200 42950 13252 43002
rect 4376 42406 4428 42458
rect 4440 42406 4492 42458
rect 4504 42406 4556 42458
rect 4568 42406 4620 42458
rect 4632 42406 4684 42458
rect 7803 42406 7855 42458
rect 7867 42406 7919 42458
rect 7931 42406 7983 42458
rect 7995 42406 8047 42458
rect 8059 42406 8111 42458
rect 11230 42406 11282 42458
rect 11294 42406 11346 42458
rect 11358 42406 11410 42458
rect 11422 42406 11474 42458
rect 11486 42406 11538 42458
rect 14657 42406 14709 42458
rect 14721 42406 14773 42458
rect 14785 42406 14837 42458
rect 14849 42406 14901 42458
rect 14913 42406 14965 42458
rect 2663 41862 2715 41914
rect 2727 41862 2779 41914
rect 2791 41862 2843 41914
rect 2855 41862 2907 41914
rect 2919 41862 2971 41914
rect 6090 41862 6142 41914
rect 6154 41862 6206 41914
rect 6218 41862 6270 41914
rect 6282 41862 6334 41914
rect 6346 41862 6398 41914
rect 9517 41862 9569 41914
rect 9581 41862 9633 41914
rect 9645 41862 9697 41914
rect 9709 41862 9761 41914
rect 9773 41862 9825 41914
rect 12944 41862 12996 41914
rect 13008 41862 13060 41914
rect 13072 41862 13124 41914
rect 13136 41862 13188 41914
rect 13200 41862 13252 41914
rect 4376 41318 4428 41370
rect 4440 41318 4492 41370
rect 4504 41318 4556 41370
rect 4568 41318 4620 41370
rect 4632 41318 4684 41370
rect 7803 41318 7855 41370
rect 7867 41318 7919 41370
rect 7931 41318 7983 41370
rect 7995 41318 8047 41370
rect 8059 41318 8111 41370
rect 11230 41318 11282 41370
rect 11294 41318 11346 41370
rect 11358 41318 11410 41370
rect 11422 41318 11474 41370
rect 11486 41318 11538 41370
rect 14657 41318 14709 41370
rect 14721 41318 14773 41370
rect 14785 41318 14837 41370
rect 14849 41318 14901 41370
rect 14913 41318 14965 41370
rect 2663 40774 2715 40826
rect 2727 40774 2779 40826
rect 2791 40774 2843 40826
rect 2855 40774 2907 40826
rect 2919 40774 2971 40826
rect 6090 40774 6142 40826
rect 6154 40774 6206 40826
rect 6218 40774 6270 40826
rect 6282 40774 6334 40826
rect 6346 40774 6398 40826
rect 9517 40774 9569 40826
rect 9581 40774 9633 40826
rect 9645 40774 9697 40826
rect 9709 40774 9761 40826
rect 9773 40774 9825 40826
rect 12944 40774 12996 40826
rect 13008 40774 13060 40826
rect 13072 40774 13124 40826
rect 13136 40774 13188 40826
rect 13200 40774 13252 40826
rect 4376 40230 4428 40282
rect 4440 40230 4492 40282
rect 4504 40230 4556 40282
rect 4568 40230 4620 40282
rect 4632 40230 4684 40282
rect 7803 40230 7855 40282
rect 7867 40230 7919 40282
rect 7931 40230 7983 40282
rect 7995 40230 8047 40282
rect 8059 40230 8111 40282
rect 11230 40230 11282 40282
rect 11294 40230 11346 40282
rect 11358 40230 11410 40282
rect 11422 40230 11474 40282
rect 11486 40230 11538 40282
rect 14657 40230 14709 40282
rect 14721 40230 14773 40282
rect 14785 40230 14837 40282
rect 14849 40230 14901 40282
rect 14913 40230 14965 40282
rect 2663 39686 2715 39738
rect 2727 39686 2779 39738
rect 2791 39686 2843 39738
rect 2855 39686 2907 39738
rect 2919 39686 2971 39738
rect 6090 39686 6142 39738
rect 6154 39686 6206 39738
rect 6218 39686 6270 39738
rect 6282 39686 6334 39738
rect 6346 39686 6398 39738
rect 9517 39686 9569 39738
rect 9581 39686 9633 39738
rect 9645 39686 9697 39738
rect 9709 39686 9761 39738
rect 9773 39686 9825 39738
rect 12944 39686 12996 39738
rect 13008 39686 13060 39738
rect 13072 39686 13124 39738
rect 13136 39686 13188 39738
rect 13200 39686 13252 39738
rect 4376 39142 4428 39194
rect 4440 39142 4492 39194
rect 4504 39142 4556 39194
rect 4568 39142 4620 39194
rect 4632 39142 4684 39194
rect 7803 39142 7855 39194
rect 7867 39142 7919 39194
rect 7931 39142 7983 39194
rect 7995 39142 8047 39194
rect 8059 39142 8111 39194
rect 11230 39142 11282 39194
rect 11294 39142 11346 39194
rect 11358 39142 11410 39194
rect 11422 39142 11474 39194
rect 11486 39142 11538 39194
rect 14657 39142 14709 39194
rect 14721 39142 14773 39194
rect 14785 39142 14837 39194
rect 14849 39142 14901 39194
rect 14913 39142 14965 39194
rect 2663 38598 2715 38650
rect 2727 38598 2779 38650
rect 2791 38598 2843 38650
rect 2855 38598 2907 38650
rect 2919 38598 2971 38650
rect 6090 38598 6142 38650
rect 6154 38598 6206 38650
rect 6218 38598 6270 38650
rect 6282 38598 6334 38650
rect 6346 38598 6398 38650
rect 9517 38598 9569 38650
rect 9581 38598 9633 38650
rect 9645 38598 9697 38650
rect 9709 38598 9761 38650
rect 9773 38598 9825 38650
rect 12944 38598 12996 38650
rect 13008 38598 13060 38650
rect 13072 38598 13124 38650
rect 13136 38598 13188 38650
rect 13200 38598 13252 38650
rect 4376 38054 4428 38106
rect 4440 38054 4492 38106
rect 4504 38054 4556 38106
rect 4568 38054 4620 38106
rect 4632 38054 4684 38106
rect 7803 38054 7855 38106
rect 7867 38054 7919 38106
rect 7931 38054 7983 38106
rect 7995 38054 8047 38106
rect 8059 38054 8111 38106
rect 11230 38054 11282 38106
rect 11294 38054 11346 38106
rect 11358 38054 11410 38106
rect 11422 38054 11474 38106
rect 11486 38054 11538 38106
rect 14657 38054 14709 38106
rect 14721 38054 14773 38106
rect 14785 38054 14837 38106
rect 14849 38054 14901 38106
rect 14913 38054 14965 38106
rect 2663 37510 2715 37562
rect 2727 37510 2779 37562
rect 2791 37510 2843 37562
rect 2855 37510 2907 37562
rect 2919 37510 2971 37562
rect 6090 37510 6142 37562
rect 6154 37510 6206 37562
rect 6218 37510 6270 37562
rect 6282 37510 6334 37562
rect 6346 37510 6398 37562
rect 9517 37510 9569 37562
rect 9581 37510 9633 37562
rect 9645 37510 9697 37562
rect 9709 37510 9761 37562
rect 9773 37510 9825 37562
rect 12944 37510 12996 37562
rect 13008 37510 13060 37562
rect 13072 37510 13124 37562
rect 13136 37510 13188 37562
rect 13200 37510 13252 37562
rect 4376 36966 4428 37018
rect 4440 36966 4492 37018
rect 4504 36966 4556 37018
rect 4568 36966 4620 37018
rect 4632 36966 4684 37018
rect 7803 36966 7855 37018
rect 7867 36966 7919 37018
rect 7931 36966 7983 37018
rect 7995 36966 8047 37018
rect 8059 36966 8111 37018
rect 11230 36966 11282 37018
rect 11294 36966 11346 37018
rect 11358 36966 11410 37018
rect 11422 36966 11474 37018
rect 11486 36966 11538 37018
rect 14657 36966 14709 37018
rect 14721 36966 14773 37018
rect 14785 36966 14837 37018
rect 14849 36966 14901 37018
rect 14913 36966 14965 37018
rect 2663 36422 2715 36474
rect 2727 36422 2779 36474
rect 2791 36422 2843 36474
rect 2855 36422 2907 36474
rect 2919 36422 2971 36474
rect 6090 36422 6142 36474
rect 6154 36422 6206 36474
rect 6218 36422 6270 36474
rect 6282 36422 6334 36474
rect 6346 36422 6398 36474
rect 9517 36422 9569 36474
rect 9581 36422 9633 36474
rect 9645 36422 9697 36474
rect 9709 36422 9761 36474
rect 9773 36422 9825 36474
rect 12944 36422 12996 36474
rect 13008 36422 13060 36474
rect 13072 36422 13124 36474
rect 13136 36422 13188 36474
rect 13200 36422 13252 36474
rect 14464 36023 14516 36032
rect 14464 35989 14473 36023
rect 14473 35989 14507 36023
rect 14507 35989 14516 36023
rect 14464 35980 14516 35989
rect 4376 35878 4428 35930
rect 4440 35878 4492 35930
rect 4504 35878 4556 35930
rect 4568 35878 4620 35930
rect 4632 35878 4684 35930
rect 7803 35878 7855 35930
rect 7867 35878 7919 35930
rect 7931 35878 7983 35930
rect 7995 35878 8047 35930
rect 8059 35878 8111 35930
rect 11230 35878 11282 35930
rect 11294 35878 11346 35930
rect 11358 35878 11410 35930
rect 11422 35878 11474 35930
rect 11486 35878 11538 35930
rect 14657 35878 14709 35930
rect 14721 35878 14773 35930
rect 14785 35878 14837 35930
rect 14849 35878 14901 35930
rect 14913 35878 14965 35930
rect 2663 35334 2715 35386
rect 2727 35334 2779 35386
rect 2791 35334 2843 35386
rect 2855 35334 2907 35386
rect 2919 35334 2971 35386
rect 6090 35334 6142 35386
rect 6154 35334 6206 35386
rect 6218 35334 6270 35386
rect 6282 35334 6334 35386
rect 6346 35334 6398 35386
rect 9517 35334 9569 35386
rect 9581 35334 9633 35386
rect 9645 35334 9697 35386
rect 9709 35334 9761 35386
rect 9773 35334 9825 35386
rect 12944 35334 12996 35386
rect 13008 35334 13060 35386
rect 13072 35334 13124 35386
rect 13136 35334 13188 35386
rect 13200 35334 13252 35386
rect 4376 34790 4428 34842
rect 4440 34790 4492 34842
rect 4504 34790 4556 34842
rect 4568 34790 4620 34842
rect 4632 34790 4684 34842
rect 7803 34790 7855 34842
rect 7867 34790 7919 34842
rect 7931 34790 7983 34842
rect 7995 34790 8047 34842
rect 8059 34790 8111 34842
rect 11230 34790 11282 34842
rect 11294 34790 11346 34842
rect 11358 34790 11410 34842
rect 11422 34790 11474 34842
rect 11486 34790 11538 34842
rect 14657 34790 14709 34842
rect 14721 34790 14773 34842
rect 14785 34790 14837 34842
rect 14849 34790 14901 34842
rect 14913 34790 14965 34842
rect 2663 34246 2715 34298
rect 2727 34246 2779 34298
rect 2791 34246 2843 34298
rect 2855 34246 2907 34298
rect 2919 34246 2971 34298
rect 6090 34246 6142 34298
rect 6154 34246 6206 34298
rect 6218 34246 6270 34298
rect 6282 34246 6334 34298
rect 6346 34246 6398 34298
rect 9517 34246 9569 34298
rect 9581 34246 9633 34298
rect 9645 34246 9697 34298
rect 9709 34246 9761 34298
rect 9773 34246 9825 34298
rect 12944 34246 12996 34298
rect 13008 34246 13060 34298
rect 13072 34246 13124 34298
rect 13136 34246 13188 34298
rect 13200 34246 13252 34298
rect 4376 33702 4428 33754
rect 4440 33702 4492 33754
rect 4504 33702 4556 33754
rect 4568 33702 4620 33754
rect 4632 33702 4684 33754
rect 7803 33702 7855 33754
rect 7867 33702 7919 33754
rect 7931 33702 7983 33754
rect 7995 33702 8047 33754
rect 8059 33702 8111 33754
rect 11230 33702 11282 33754
rect 11294 33702 11346 33754
rect 11358 33702 11410 33754
rect 11422 33702 11474 33754
rect 11486 33702 11538 33754
rect 14657 33702 14709 33754
rect 14721 33702 14773 33754
rect 14785 33702 14837 33754
rect 14849 33702 14901 33754
rect 14913 33702 14965 33754
rect 2663 33158 2715 33210
rect 2727 33158 2779 33210
rect 2791 33158 2843 33210
rect 2855 33158 2907 33210
rect 2919 33158 2971 33210
rect 6090 33158 6142 33210
rect 6154 33158 6206 33210
rect 6218 33158 6270 33210
rect 6282 33158 6334 33210
rect 6346 33158 6398 33210
rect 9517 33158 9569 33210
rect 9581 33158 9633 33210
rect 9645 33158 9697 33210
rect 9709 33158 9761 33210
rect 9773 33158 9825 33210
rect 12944 33158 12996 33210
rect 13008 33158 13060 33210
rect 13072 33158 13124 33210
rect 13136 33158 13188 33210
rect 13200 33158 13252 33210
rect 4376 32614 4428 32666
rect 4440 32614 4492 32666
rect 4504 32614 4556 32666
rect 4568 32614 4620 32666
rect 4632 32614 4684 32666
rect 7803 32614 7855 32666
rect 7867 32614 7919 32666
rect 7931 32614 7983 32666
rect 7995 32614 8047 32666
rect 8059 32614 8111 32666
rect 11230 32614 11282 32666
rect 11294 32614 11346 32666
rect 11358 32614 11410 32666
rect 11422 32614 11474 32666
rect 11486 32614 11538 32666
rect 14657 32614 14709 32666
rect 14721 32614 14773 32666
rect 14785 32614 14837 32666
rect 14849 32614 14901 32666
rect 14913 32614 14965 32666
rect 2663 32070 2715 32122
rect 2727 32070 2779 32122
rect 2791 32070 2843 32122
rect 2855 32070 2907 32122
rect 2919 32070 2971 32122
rect 6090 32070 6142 32122
rect 6154 32070 6206 32122
rect 6218 32070 6270 32122
rect 6282 32070 6334 32122
rect 6346 32070 6398 32122
rect 9517 32070 9569 32122
rect 9581 32070 9633 32122
rect 9645 32070 9697 32122
rect 9709 32070 9761 32122
rect 9773 32070 9825 32122
rect 12944 32070 12996 32122
rect 13008 32070 13060 32122
rect 13072 32070 13124 32122
rect 13136 32070 13188 32122
rect 13200 32070 13252 32122
rect 4376 31526 4428 31578
rect 4440 31526 4492 31578
rect 4504 31526 4556 31578
rect 4568 31526 4620 31578
rect 4632 31526 4684 31578
rect 7803 31526 7855 31578
rect 7867 31526 7919 31578
rect 7931 31526 7983 31578
rect 7995 31526 8047 31578
rect 8059 31526 8111 31578
rect 11230 31526 11282 31578
rect 11294 31526 11346 31578
rect 11358 31526 11410 31578
rect 11422 31526 11474 31578
rect 11486 31526 11538 31578
rect 14657 31526 14709 31578
rect 14721 31526 14773 31578
rect 14785 31526 14837 31578
rect 14849 31526 14901 31578
rect 14913 31526 14965 31578
rect 2663 30982 2715 31034
rect 2727 30982 2779 31034
rect 2791 30982 2843 31034
rect 2855 30982 2907 31034
rect 2919 30982 2971 31034
rect 6090 30982 6142 31034
rect 6154 30982 6206 31034
rect 6218 30982 6270 31034
rect 6282 30982 6334 31034
rect 6346 30982 6398 31034
rect 9517 30982 9569 31034
rect 9581 30982 9633 31034
rect 9645 30982 9697 31034
rect 9709 30982 9761 31034
rect 9773 30982 9825 31034
rect 12944 30982 12996 31034
rect 13008 30982 13060 31034
rect 13072 30982 13124 31034
rect 13136 30982 13188 31034
rect 13200 30982 13252 31034
rect 4376 30438 4428 30490
rect 4440 30438 4492 30490
rect 4504 30438 4556 30490
rect 4568 30438 4620 30490
rect 4632 30438 4684 30490
rect 7803 30438 7855 30490
rect 7867 30438 7919 30490
rect 7931 30438 7983 30490
rect 7995 30438 8047 30490
rect 8059 30438 8111 30490
rect 11230 30438 11282 30490
rect 11294 30438 11346 30490
rect 11358 30438 11410 30490
rect 11422 30438 11474 30490
rect 11486 30438 11538 30490
rect 14657 30438 14709 30490
rect 14721 30438 14773 30490
rect 14785 30438 14837 30490
rect 14849 30438 14901 30490
rect 14913 30438 14965 30490
rect 2663 29894 2715 29946
rect 2727 29894 2779 29946
rect 2791 29894 2843 29946
rect 2855 29894 2907 29946
rect 2919 29894 2971 29946
rect 6090 29894 6142 29946
rect 6154 29894 6206 29946
rect 6218 29894 6270 29946
rect 6282 29894 6334 29946
rect 6346 29894 6398 29946
rect 9517 29894 9569 29946
rect 9581 29894 9633 29946
rect 9645 29894 9697 29946
rect 9709 29894 9761 29946
rect 9773 29894 9825 29946
rect 12944 29894 12996 29946
rect 13008 29894 13060 29946
rect 13072 29894 13124 29946
rect 13136 29894 13188 29946
rect 13200 29894 13252 29946
rect 4376 29350 4428 29402
rect 4440 29350 4492 29402
rect 4504 29350 4556 29402
rect 4568 29350 4620 29402
rect 4632 29350 4684 29402
rect 7803 29350 7855 29402
rect 7867 29350 7919 29402
rect 7931 29350 7983 29402
rect 7995 29350 8047 29402
rect 8059 29350 8111 29402
rect 11230 29350 11282 29402
rect 11294 29350 11346 29402
rect 11358 29350 11410 29402
rect 11422 29350 11474 29402
rect 11486 29350 11538 29402
rect 14657 29350 14709 29402
rect 14721 29350 14773 29402
rect 14785 29350 14837 29402
rect 14849 29350 14901 29402
rect 14913 29350 14965 29402
rect 2663 28806 2715 28858
rect 2727 28806 2779 28858
rect 2791 28806 2843 28858
rect 2855 28806 2907 28858
rect 2919 28806 2971 28858
rect 6090 28806 6142 28858
rect 6154 28806 6206 28858
rect 6218 28806 6270 28858
rect 6282 28806 6334 28858
rect 6346 28806 6398 28858
rect 9517 28806 9569 28858
rect 9581 28806 9633 28858
rect 9645 28806 9697 28858
rect 9709 28806 9761 28858
rect 9773 28806 9825 28858
rect 12944 28806 12996 28858
rect 13008 28806 13060 28858
rect 13072 28806 13124 28858
rect 13136 28806 13188 28858
rect 13200 28806 13252 28858
rect 4376 28262 4428 28314
rect 4440 28262 4492 28314
rect 4504 28262 4556 28314
rect 4568 28262 4620 28314
rect 4632 28262 4684 28314
rect 7803 28262 7855 28314
rect 7867 28262 7919 28314
rect 7931 28262 7983 28314
rect 7995 28262 8047 28314
rect 8059 28262 8111 28314
rect 11230 28262 11282 28314
rect 11294 28262 11346 28314
rect 11358 28262 11410 28314
rect 11422 28262 11474 28314
rect 11486 28262 11538 28314
rect 14657 28262 14709 28314
rect 14721 28262 14773 28314
rect 14785 28262 14837 28314
rect 14849 28262 14901 28314
rect 14913 28262 14965 28314
rect 14464 27999 14516 28008
rect 14464 27965 14473 27999
rect 14473 27965 14507 27999
rect 14507 27965 14516 27999
rect 14464 27956 14516 27965
rect 2663 27718 2715 27770
rect 2727 27718 2779 27770
rect 2791 27718 2843 27770
rect 2855 27718 2907 27770
rect 2919 27718 2971 27770
rect 6090 27718 6142 27770
rect 6154 27718 6206 27770
rect 6218 27718 6270 27770
rect 6282 27718 6334 27770
rect 6346 27718 6398 27770
rect 9517 27718 9569 27770
rect 9581 27718 9633 27770
rect 9645 27718 9697 27770
rect 9709 27718 9761 27770
rect 9773 27718 9825 27770
rect 12944 27718 12996 27770
rect 13008 27718 13060 27770
rect 13072 27718 13124 27770
rect 13136 27718 13188 27770
rect 13200 27718 13252 27770
rect 4376 27174 4428 27226
rect 4440 27174 4492 27226
rect 4504 27174 4556 27226
rect 4568 27174 4620 27226
rect 4632 27174 4684 27226
rect 7803 27174 7855 27226
rect 7867 27174 7919 27226
rect 7931 27174 7983 27226
rect 7995 27174 8047 27226
rect 8059 27174 8111 27226
rect 11230 27174 11282 27226
rect 11294 27174 11346 27226
rect 11358 27174 11410 27226
rect 11422 27174 11474 27226
rect 11486 27174 11538 27226
rect 14657 27174 14709 27226
rect 14721 27174 14773 27226
rect 14785 27174 14837 27226
rect 14849 27174 14901 27226
rect 14913 27174 14965 27226
rect 2663 26630 2715 26682
rect 2727 26630 2779 26682
rect 2791 26630 2843 26682
rect 2855 26630 2907 26682
rect 2919 26630 2971 26682
rect 6090 26630 6142 26682
rect 6154 26630 6206 26682
rect 6218 26630 6270 26682
rect 6282 26630 6334 26682
rect 6346 26630 6398 26682
rect 9517 26630 9569 26682
rect 9581 26630 9633 26682
rect 9645 26630 9697 26682
rect 9709 26630 9761 26682
rect 9773 26630 9825 26682
rect 12944 26630 12996 26682
rect 13008 26630 13060 26682
rect 13072 26630 13124 26682
rect 13136 26630 13188 26682
rect 13200 26630 13252 26682
rect 4376 26086 4428 26138
rect 4440 26086 4492 26138
rect 4504 26086 4556 26138
rect 4568 26086 4620 26138
rect 4632 26086 4684 26138
rect 7803 26086 7855 26138
rect 7867 26086 7919 26138
rect 7931 26086 7983 26138
rect 7995 26086 8047 26138
rect 8059 26086 8111 26138
rect 11230 26086 11282 26138
rect 11294 26086 11346 26138
rect 11358 26086 11410 26138
rect 11422 26086 11474 26138
rect 11486 26086 11538 26138
rect 14657 26086 14709 26138
rect 14721 26086 14773 26138
rect 14785 26086 14837 26138
rect 14849 26086 14901 26138
rect 14913 26086 14965 26138
rect 2663 25542 2715 25594
rect 2727 25542 2779 25594
rect 2791 25542 2843 25594
rect 2855 25542 2907 25594
rect 2919 25542 2971 25594
rect 6090 25542 6142 25594
rect 6154 25542 6206 25594
rect 6218 25542 6270 25594
rect 6282 25542 6334 25594
rect 6346 25542 6398 25594
rect 9517 25542 9569 25594
rect 9581 25542 9633 25594
rect 9645 25542 9697 25594
rect 9709 25542 9761 25594
rect 9773 25542 9825 25594
rect 12944 25542 12996 25594
rect 13008 25542 13060 25594
rect 13072 25542 13124 25594
rect 13136 25542 13188 25594
rect 13200 25542 13252 25594
rect 4376 24998 4428 25050
rect 4440 24998 4492 25050
rect 4504 24998 4556 25050
rect 4568 24998 4620 25050
rect 4632 24998 4684 25050
rect 7803 24998 7855 25050
rect 7867 24998 7919 25050
rect 7931 24998 7983 25050
rect 7995 24998 8047 25050
rect 8059 24998 8111 25050
rect 11230 24998 11282 25050
rect 11294 24998 11346 25050
rect 11358 24998 11410 25050
rect 11422 24998 11474 25050
rect 11486 24998 11538 25050
rect 14657 24998 14709 25050
rect 14721 24998 14773 25050
rect 14785 24998 14837 25050
rect 14849 24998 14901 25050
rect 14913 24998 14965 25050
rect 2663 24454 2715 24506
rect 2727 24454 2779 24506
rect 2791 24454 2843 24506
rect 2855 24454 2907 24506
rect 2919 24454 2971 24506
rect 6090 24454 6142 24506
rect 6154 24454 6206 24506
rect 6218 24454 6270 24506
rect 6282 24454 6334 24506
rect 6346 24454 6398 24506
rect 9517 24454 9569 24506
rect 9581 24454 9633 24506
rect 9645 24454 9697 24506
rect 9709 24454 9761 24506
rect 9773 24454 9825 24506
rect 12944 24454 12996 24506
rect 13008 24454 13060 24506
rect 13072 24454 13124 24506
rect 13136 24454 13188 24506
rect 13200 24454 13252 24506
rect 4376 23910 4428 23962
rect 4440 23910 4492 23962
rect 4504 23910 4556 23962
rect 4568 23910 4620 23962
rect 4632 23910 4684 23962
rect 7803 23910 7855 23962
rect 7867 23910 7919 23962
rect 7931 23910 7983 23962
rect 7995 23910 8047 23962
rect 8059 23910 8111 23962
rect 11230 23910 11282 23962
rect 11294 23910 11346 23962
rect 11358 23910 11410 23962
rect 11422 23910 11474 23962
rect 11486 23910 11538 23962
rect 14657 23910 14709 23962
rect 14721 23910 14773 23962
rect 14785 23910 14837 23962
rect 14849 23910 14901 23962
rect 14913 23910 14965 23962
rect 2663 23366 2715 23418
rect 2727 23366 2779 23418
rect 2791 23366 2843 23418
rect 2855 23366 2907 23418
rect 2919 23366 2971 23418
rect 6090 23366 6142 23418
rect 6154 23366 6206 23418
rect 6218 23366 6270 23418
rect 6282 23366 6334 23418
rect 6346 23366 6398 23418
rect 9517 23366 9569 23418
rect 9581 23366 9633 23418
rect 9645 23366 9697 23418
rect 9709 23366 9761 23418
rect 9773 23366 9825 23418
rect 12944 23366 12996 23418
rect 13008 23366 13060 23418
rect 13072 23366 13124 23418
rect 13136 23366 13188 23418
rect 13200 23366 13252 23418
rect 4376 22822 4428 22874
rect 4440 22822 4492 22874
rect 4504 22822 4556 22874
rect 4568 22822 4620 22874
rect 4632 22822 4684 22874
rect 7803 22822 7855 22874
rect 7867 22822 7919 22874
rect 7931 22822 7983 22874
rect 7995 22822 8047 22874
rect 8059 22822 8111 22874
rect 11230 22822 11282 22874
rect 11294 22822 11346 22874
rect 11358 22822 11410 22874
rect 11422 22822 11474 22874
rect 11486 22822 11538 22874
rect 14657 22822 14709 22874
rect 14721 22822 14773 22874
rect 14785 22822 14837 22874
rect 14849 22822 14901 22874
rect 14913 22822 14965 22874
rect 2663 22278 2715 22330
rect 2727 22278 2779 22330
rect 2791 22278 2843 22330
rect 2855 22278 2907 22330
rect 2919 22278 2971 22330
rect 6090 22278 6142 22330
rect 6154 22278 6206 22330
rect 6218 22278 6270 22330
rect 6282 22278 6334 22330
rect 6346 22278 6398 22330
rect 9517 22278 9569 22330
rect 9581 22278 9633 22330
rect 9645 22278 9697 22330
rect 9709 22278 9761 22330
rect 9773 22278 9825 22330
rect 12944 22278 12996 22330
rect 13008 22278 13060 22330
rect 13072 22278 13124 22330
rect 13136 22278 13188 22330
rect 13200 22278 13252 22330
rect 4376 21734 4428 21786
rect 4440 21734 4492 21786
rect 4504 21734 4556 21786
rect 4568 21734 4620 21786
rect 4632 21734 4684 21786
rect 7803 21734 7855 21786
rect 7867 21734 7919 21786
rect 7931 21734 7983 21786
rect 7995 21734 8047 21786
rect 8059 21734 8111 21786
rect 11230 21734 11282 21786
rect 11294 21734 11346 21786
rect 11358 21734 11410 21786
rect 11422 21734 11474 21786
rect 11486 21734 11538 21786
rect 14657 21734 14709 21786
rect 14721 21734 14773 21786
rect 14785 21734 14837 21786
rect 14849 21734 14901 21786
rect 14913 21734 14965 21786
rect 2663 21190 2715 21242
rect 2727 21190 2779 21242
rect 2791 21190 2843 21242
rect 2855 21190 2907 21242
rect 2919 21190 2971 21242
rect 6090 21190 6142 21242
rect 6154 21190 6206 21242
rect 6218 21190 6270 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 9517 21190 9569 21242
rect 9581 21190 9633 21242
rect 9645 21190 9697 21242
rect 9709 21190 9761 21242
rect 9773 21190 9825 21242
rect 12944 21190 12996 21242
rect 13008 21190 13060 21242
rect 13072 21190 13124 21242
rect 13136 21190 13188 21242
rect 13200 21190 13252 21242
rect 4376 20646 4428 20698
rect 4440 20646 4492 20698
rect 4504 20646 4556 20698
rect 4568 20646 4620 20698
rect 4632 20646 4684 20698
rect 7803 20646 7855 20698
rect 7867 20646 7919 20698
rect 7931 20646 7983 20698
rect 7995 20646 8047 20698
rect 8059 20646 8111 20698
rect 11230 20646 11282 20698
rect 11294 20646 11346 20698
rect 11358 20646 11410 20698
rect 11422 20646 11474 20698
rect 11486 20646 11538 20698
rect 14657 20646 14709 20698
rect 14721 20646 14773 20698
rect 14785 20646 14837 20698
rect 14849 20646 14901 20698
rect 14913 20646 14965 20698
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 2663 20102 2715 20154
rect 2727 20102 2779 20154
rect 2791 20102 2843 20154
rect 2855 20102 2907 20154
rect 2919 20102 2971 20154
rect 6090 20102 6142 20154
rect 6154 20102 6206 20154
rect 6218 20102 6270 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 9517 20102 9569 20154
rect 9581 20102 9633 20154
rect 9645 20102 9697 20154
rect 9709 20102 9761 20154
rect 9773 20102 9825 20154
rect 12944 20102 12996 20154
rect 13008 20102 13060 20154
rect 13072 20102 13124 20154
rect 13136 20102 13188 20154
rect 13200 20102 13252 20154
rect 4376 19558 4428 19610
rect 4440 19558 4492 19610
rect 4504 19558 4556 19610
rect 4568 19558 4620 19610
rect 4632 19558 4684 19610
rect 7803 19558 7855 19610
rect 7867 19558 7919 19610
rect 7931 19558 7983 19610
rect 7995 19558 8047 19610
rect 8059 19558 8111 19610
rect 11230 19558 11282 19610
rect 11294 19558 11346 19610
rect 11358 19558 11410 19610
rect 11422 19558 11474 19610
rect 11486 19558 11538 19610
rect 14657 19558 14709 19610
rect 14721 19558 14773 19610
rect 14785 19558 14837 19610
rect 14849 19558 14901 19610
rect 14913 19558 14965 19610
rect 2663 19014 2715 19066
rect 2727 19014 2779 19066
rect 2791 19014 2843 19066
rect 2855 19014 2907 19066
rect 2919 19014 2971 19066
rect 6090 19014 6142 19066
rect 6154 19014 6206 19066
rect 6218 19014 6270 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 9517 19014 9569 19066
rect 9581 19014 9633 19066
rect 9645 19014 9697 19066
rect 9709 19014 9761 19066
rect 9773 19014 9825 19066
rect 12944 19014 12996 19066
rect 13008 19014 13060 19066
rect 13072 19014 13124 19066
rect 13136 19014 13188 19066
rect 13200 19014 13252 19066
rect 4376 18470 4428 18522
rect 4440 18470 4492 18522
rect 4504 18470 4556 18522
rect 4568 18470 4620 18522
rect 4632 18470 4684 18522
rect 7803 18470 7855 18522
rect 7867 18470 7919 18522
rect 7931 18470 7983 18522
rect 7995 18470 8047 18522
rect 8059 18470 8111 18522
rect 11230 18470 11282 18522
rect 11294 18470 11346 18522
rect 11358 18470 11410 18522
rect 11422 18470 11474 18522
rect 11486 18470 11538 18522
rect 14657 18470 14709 18522
rect 14721 18470 14773 18522
rect 14785 18470 14837 18522
rect 14849 18470 14901 18522
rect 14913 18470 14965 18522
rect 2663 17926 2715 17978
rect 2727 17926 2779 17978
rect 2791 17926 2843 17978
rect 2855 17926 2907 17978
rect 2919 17926 2971 17978
rect 6090 17926 6142 17978
rect 6154 17926 6206 17978
rect 6218 17926 6270 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 9517 17926 9569 17978
rect 9581 17926 9633 17978
rect 9645 17926 9697 17978
rect 9709 17926 9761 17978
rect 9773 17926 9825 17978
rect 12944 17926 12996 17978
rect 13008 17926 13060 17978
rect 13072 17926 13124 17978
rect 13136 17926 13188 17978
rect 13200 17926 13252 17978
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 14464 12155 14516 12164
rect 14464 12121 14473 12155
rect 14473 12121 14507 12155
rect 14507 12121 14516 12155
rect 14464 12112 14516 12121
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
<< metal2 >>
rect 4376 45724 4684 45733
rect 4376 45722 4382 45724
rect 4438 45722 4462 45724
rect 4518 45722 4542 45724
rect 4598 45722 4622 45724
rect 4678 45722 4684 45724
rect 4438 45670 4440 45722
rect 4620 45670 4622 45722
rect 4376 45668 4382 45670
rect 4438 45668 4462 45670
rect 4518 45668 4542 45670
rect 4598 45668 4622 45670
rect 4678 45668 4684 45670
rect 4376 45659 4684 45668
rect 7803 45724 8111 45733
rect 7803 45722 7809 45724
rect 7865 45722 7889 45724
rect 7945 45722 7969 45724
rect 8025 45722 8049 45724
rect 8105 45722 8111 45724
rect 7865 45670 7867 45722
rect 8047 45670 8049 45722
rect 7803 45668 7809 45670
rect 7865 45668 7889 45670
rect 7945 45668 7969 45670
rect 8025 45668 8049 45670
rect 8105 45668 8111 45670
rect 7803 45659 8111 45668
rect 11230 45724 11538 45733
rect 11230 45722 11236 45724
rect 11292 45722 11316 45724
rect 11372 45722 11396 45724
rect 11452 45722 11476 45724
rect 11532 45722 11538 45724
rect 11292 45670 11294 45722
rect 11474 45670 11476 45722
rect 11230 45668 11236 45670
rect 11292 45668 11316 45670
rect 11372 45668 11396 45670
rect 11452 45668 11476 45670
rect 11532 45668 11538 45670
rect 11230 45659 11538 45668
rect 14657 45724 14965 45733
rect 14657 45722 14663 45724
rect 14719 45722 14743 45724
rect 14799 45722 14823 45724
rect 14879 45722 14903 45724
rect 14959 45722 14965 45724
rect 14719 45670 14721 45722
rect 14901 45670 14903 45722
rect 14657 45668 14663 45670
rect 14719 45668 14743 45670
rect 14799 45668 14823 45670
rect 14879 45668 14903 45670
rect 14959 45668 14965 45670
rect 14657 45659 14965 45668
rect 2663 45180 2971 45189
rect 2663 45178 2669 45180
rect 2725 45178 2749 45180
rect 2805 45178 2829 45180
rect 2885 45178 2909 45180
rect 2965 45178 2971 45180
rect 2725 45126 2727 45178
rect 2907 45126 2909 45178
rect 2663 45124 2669 45126
rect 2725 45124 2749 45126
rect 2805 45124 2829 45126
rect 2885 45124 2909 45126
rect 2965 45124 2971 45126
rect 2663 45115 2971 45124
rect 6090 45180 6398 45189
rect 6090 45178 6096 45180
rect 6152 45178 6176 45180
rect 6232 45178 6256 45180
rect 6312 45178 6336 45180
rect 6392 45178 6398 45180
rect 6152 45126 6154 45178
rect 6334 45126 6336 45178
rect 6090 45124 6096 45126
rect 6152 45124 6176 45126
rect 6232 45124 6256 45126
rect 6312 45124 6336 45126
rect 6392 45124 6398 45126
rect 6090 45115 6398 45124
rect 9517 45180 9825 45189
rect 9517 45178 9523 45180
rect 9579 45178 9603 45180
rect 9659 45178 9683 45180
rect 9739 45178 9763 45180
rect 9819 45178 9825 45180
rect 9579 45126 9581 45178
rect 9761 45126 9763 45178
rect 9517 45124 9523 45126
rect 9579 45124 9603 45126
rect 9659 45124 9683 45126
rect 9739 45124 9763 45126
rect 9819 45124 9825 45126
rect 9517 45115 9825 45124
rect 12944 45180 13252 45189
rect 12944 45178 12950 45180
rect 13006 45178 13030 45180
rect 13086 45178 13110 45180
rect 13166 45178 13190 45180
rect 13246 45178 13252 45180
rect 13006 45126 13008 45178
rect 13188 45126 13190 45178
rect 12944 45124 12950 45126
rect 13006 45124 13030 45126
rect 13086 45124 13110 45126
rect 13166 45124 13190 45126
rect 13246 45124 13252 45126
rect 12944 45115 13252 45124
rect 4376 44636 4684 44645
rect 4376 44634 4382 44636
rect 4438 44634 4462 44636
rect 4518 44634 4542 44636
rect 4598 44634 4622 44636
rect 4678 44634 4684 44636
rect 4438 44582 4440 44634
rect 4620 44582 4622 44634
rect 4376 44580 4382 44582
rect 4438 44580 4462 44582
rect 4518 44580 4542 44582
rect 4598 44580 4622 44582
rect 4678 44580 4684 44582
rect 4376 44571 4684 44580
rect 7803 44636 8111 44645
rect 7803 44634 7809 44636
rect 7865 44634 7889 44636
rect 7945 44634 7969 44636
rect 8025 44634 8049 44636
rect 8105 44634 8111 44636
rect 7865 44582 7867 44634
rect 8047 44582 8049 44634
rect 7803 44580 7809 44582
rect 7865 44580 7889 44582
rect 7945 44580 7969 44582
rect 8025 44580 8049 44582
rect 8105 44580 8111 44582
rect 7803 44571 8111 44580
rect 11230 44636 11538 44645
rect 11230 44634 11236 44636
rect 11292 44634 11316 44636
rect 11372 44634 11396 44636
rect 11452 44634 11476 44636
rect 11532 44634 11538 44636
rect 11292 44582 11294 44634
rect 11474 44582 11476 44634
rect 11230 44580 11236 44582
rect 11292 44580 11316 44582
rect 11372 44580 11396 44582
rect 11452 44580 11476 44582
rect 11532 44580 11538 44582
rect 11230 44571 11538 44580
rect 14657 44636 14965 44645
rect 14657 44634 14663 44636
rect 14719 44634 14743 44636
rect 14799 44634 14823 44636
rect 14879 44634 14903 44636
rect 14959 44634 14965 44636
rect 14719 44582 14721 44634
rect 14901 44582 14903 44634
rect 14657 44580 14663 44582
rect 14719 44580 14743 44582
rect 14799 44580 14823 44582
rect 14879 44580 14903 44582
rect 14959 44580 14965 44582
rect 14657 44571 14965 44580
rect 2663 44092 2971 44101
rect 2663 44090 2669 44092
rect 2725 44090 2749 44092
rect 2805 44090 2829 44092
rect 2885 44090 2909 44092
rect 2965 44090 2971 44092
rect 2725 44038 2727 44090
rect 2907 44038 2909 44090
rect 2663 44036 2669 44038
rect 2725 44036 2749 44038
rect 2805 44036 2829 44038
rect 2885 44036 2909 44038
rect 2965 44036 2971 44038
rect 2663 44027 2971 44036
rect 6090 44092 6398 44101
rect 6090 44090 6096 44092
rect 6152 44090 6176 44092
rect 6232 44090 6256 44092
rect 6312 44090 6336 44092
rect 6392 44090 6398 44092
rect 6152 44038 6154 44090
rect 6334 44038 6336 44090
rect 6090 44036 6096 44038
rect 6152 44036 6176 44038
rect 6232 44036 6256 44038
rect 6312 44036 6336 44038
rect 6392 44036 6398 44038
rect 6090 44027 6398 44036
rect 9517 44092 9825 44101
rect 9517 44090 9523 44092
rect 9579 44090 9603 44092
rect 9659 44090 9683 44092
rect 9739 44090 9763 44092
rect 9819 44090 9825 44092
rect 9579 44038 9581 44090
rect 9761 44038 9763 44090
rect 9517 44036 9523 44038
rect 9579 44036 9603 44038
rect 9659 44036 9683 44038
rect 9739 44036 9763 44038
rect 9819 44036 9825 44038
rect 9517 44027 9825 44036
rect 12944 44092 13252 44101
rect 12944 44090 12950 44092
rect 13006 44090 13030 44092
rect 13086 44090 13110 44092
rect 13166 44090 13190 44092
rect 13246 44090 13252 44092
rect 13006 44038 13008 44090
rect 13188 44038 13190 44090
rect 12944 44036 12950 44038
rect 13006 44036 13030 44038
rect 13086 44036 13110 44038
rect 13166 44036 13190 44038
rect 13246 44036 13252 44038
rect 12944 44027 13252 44036
rect 14462 43752 14518 43761
rect 14462 43687 14464 43696
rect 14516 43687 14518 43696
rect 14464 43658 14516 43664
rect 4376 43548 4684 43557
rect 4376 43546 4382 43548
rect 4438 43546 4462 43548
rect 4518 43546 4542 43548
rect 4598 43546 4622 43548
rect 4678 43546 4684 43548
rect 4438 43494 4440 43546
rect 4620 43494 4622 43546
rect 4376 43492 4382 43494
rect 4438 43492 4462 43494
rect 4518 43492 4542 43494
rect 4598 43492 4622 43494
rect 4678 43492 4684 43494
rect 4376 43483 4684 43492
rect 7803 43548 8111 43557
rect 7803 43546 7809 43548
rect 7865 43546 7889 43548
rect 7945 43546 7969 43548
rect 8025 43546 8049 43548
rect 8105 43546 8111 43548
rect 7865 43494 7867 43546
rect 8047 43494 8049 43546
rect 7803 43492 7809 43494
rect 7865 43492 7889 43494
rect 7945 43492 7969 43494
rect 8025 43492 8049 43494
rect 8105 43492 8111 43494
rect 7803 43483 8111 43492
rect 11230 43548 11538 43557
rect 11230 43546 11236 43548
rect 11292 43546 11316 43548
rect 11372 43546 11396 43548
rect 11452 43546 11476 43548
rect 11532 43546 11538 43548
rect 11292 43494 11294 43546
rect 11474 43494 11476 43546
rect 11230 43492 11236 43494
rect 11292 43492 11316 43494
rect 11372 43492 11396 43494
rect 11452 43492 11476 43494
rect 11532 43492 11538 43494
rect 11230 43483 11538 43492
rect 14657 43548 14965 43557
rect 14657 43546 14663 43548
rect 14719 43546 14743 43548
rect 14799 43546 14823 43548
rect 14879 43546 14903 43548
rect 14959 43546 14965 43548
rect 14719 43494 14721 43546
rect 14901 43494 14903 43546
rect 14657 43492 14663 43494
rect 14719 43492 14743 43494
rect 14799 43492 14823 43494
rect 14879 43492 14903 43494
rect 14959 43492 14965 43494
rect 14657 43483 14965 43492
rect 2663 43004 2971 43013
rect 2663 43002 2669 43004
rect 2725 43002 2749 43004
rect 2805 43002 2829 43004
rect 2885 43002 2909 43004
rect 2965 43002 2971 43004
rect 2725 42950 2727 43002
rect 2907 42950 2909 43002
rect 2663 42948 2669 42950
rect 2725 42948 2749 42950
rect 2805 42948 2829 42950
rect 2885 42948 2909 42950
rect 2965 42948 2971 42950
rect 2663 42939 2971 42948
rect 6090 43004 6398 43013
rect 6090 43002 6096 43004
rect 6152 43002 6176 43004
rect 6232 43002 6256 43004
rect 6312 43002 6336 43004
rect 6392 43002 6398 43004
rect 6152 42950 6154 43002
rect 6334 42950 6336 43002
rect 6090 42948 6096 42950
rect 6152 42948 6176 42950
rect 6232 42948 6256 42950
rect 6312 42948 6336 42950
rect 6392 42948 6398 42950
rect 6090 42939 6398 42948
rect 9517 43004 9825 43013
rect 9517 43002 9523 43004
rect 9579 43002 9603 43004
rect 9659 43002 9683 43004
rect 9739 43002 9763 43004
rect 9819 43002 9825 43004
rect 9579 42950 9581 43002
rect 9761 42950 9763 43002
rect 9517 42948 9523 42950
rect 9579 42948 9603 42950
rect 9659 42948 9683 42950
rect 9739 42948 9763 42950
rect 9819 42948 9825 42950
rect 9517 42939 9825 42948
rect 12944 43004 13252 43013
rect 12944 43002 12950 43004
rect 13006 43002 13030 43004
rect 13086 43002 13110 43004
rect 13166 43002 13190 43004
rect 13246 43002 13252 43004
rect 13006 42950 13008 43002
rect 13188 42950 13190 43002
rect 12944 42948 12950 42950
rect 13006 42948 13030 42950
rect 13086 42948 13110 42950
rect 13166 42948 13190 42950
rect 13246 42948 13252 42950
rect 12944 42939 13252 42948
rect 4376 42460 4684 42469
rect 4376 42458 4382 42460
rect 4438 42458 4462 42460
rect 4518 42458 4542 42460
rect 4598 42458 4622 42460
rect 4678 42458 4684 42460
rect 4438 42406 4440 42458
rect 4620 42406 4622 42458
rect 4376 42404 4382 42406
rect 4438 42404 4462 42406
rect 4518 42404 4542 42406
rect 4598 42404 4622 42406
rect 4678 42404 4684 42406
rect 4376 42395 4684 42404
rect 7803 42460 8111 42469
rect 7803 42458 7809 42460
rect 7865 42458 7889 42460
rect 7945 42458 7969 42460
rect 8025 42458 8049 42460
rect 8105 42458 8111 42460
rect 7865 42406 7867 42458
rect 8047 42406 8049 42458
rect 7803 42404 7809 42406
rect 7865 42404 7889 42406
rect 7945 42404 7969 42406
rect 8025 42404 8049 42406
rect 8105 42404 8111 42406
rect 7803 42395 8111 42404
rect 11230 42460 11538 42469
rect 11230 42458 11236 42460
rect 11292 42458 11316 42460
rect 11372 42458 11396 42460
rect 11452 42458 11476 42460
rect 11532 42458 11538 42460
rect 11292 42406 11294 42458
rect 11474 42406 11476 42458
rect 11230 42404 11236 42406
rect 11292 42404 11316 42406
rect 11372 42404 11396 42406
rect 11452 42404 11476 42406
rect 11532 42404 11538 42406
rect 11230 42395 11538 42404
rect 14657 42460 14965 42469
rect 14657 42458 14663 42460
rect 14719 42458 14743 42460
rect 14799 42458 14823 42460
rect 14879 42458 14903 42460
rect 14959 42458 14965 42460
rect 14719 42406 14721 42458
rect 14901 42406 14903 42458
rect 14657 42404 14663 42406
rect 14719 42404 14743 42406
rect 14799 42404 14823 42406
rect 14879 42404 14903 42406
rect 14959 42404 14965 42406
rect 14657 42395 14965 42404
rect 2663 41916 2971 41925
rect 2663 41914 2669 41916
rect 2725 41914 2749 41916
rect 2805 41914 2829 41916
rect 2885 41914 2909 41916
rect 2965 41914 2971 41916
rect 2725 41862 2727 41914
rect 2907 41862 2909 41914
rect 2663 41860 2669 41862
rect 2725 41860 2749 41862
rect 2805 41860 2829 41862
rect 2885 41860 2909 41862
rect 2965 41860 2971 41862
rect 2663 41851 2971 41860
rect 6090 41916 6398 41925
rect 6090 41914 6096 41916
rect 6152 41914 6176 41916
rect 6232 41914 6256 41916
rect 6312 41914 6336 41916
rect 6392 41914 6398 41916
rect 6152 41862 6154 41914
rect 6334 41862 6336 41914
rect 6090 41860 6096 41862
rect 6152 41860 6176 41862
rect 6232 41860 6256 41862
rect 6312 41860 6336 41862
rect 6392 41860 6398 41862
rect 6090 41851 6398 41860
rect 9517 41916 9825 41925
rect 9517 41914 9523 41916
rect 9579 41914 9603 41916
rect 9659 41914 9683 41916
rect 9739 41914 9763 41916
rect 9819 41914 9825 41916
rect 9579 41862 9581 41914
rect 9761 41862 9763 41914
rect 9517 41860 9523 41862
rect 9579 41860 9603 41862
rect 9659 41860 9683 41862
rect 9739 41860 9763 41862
rect 9819 41860 9825 41862
rect 9517 41851 9825 41860
rect 12944 41916 13252 41925
rect 12944 41914 12950 41916
rect 13006 41914 13030 41916
rect 13086 41914 13110 41916
rect 13166 41914 13190 41916
rect 13246 41914 13252 41916
rect 13006 41862 13008 41914
rect 13188 41862 13190 41914
rect 12944 41860 12950 41862
rect 13006 41860 13030 41862
rect 13086 41860 13110 41862
rect 13166 41860 13190 41862
rect 13246 41860 13252 41862
rect 12944 41851 13252 41860
rect 4376 41372 4684 41381
rect 4376 41370 4382 41372
rect 4438 41370 4462 41372
rect 4518 41370 4542 41372
rect 4598 41370 4622 41372
rect 4678 41370 4684 41372
rect 4438 41318 4440 41370
rect 4620 41318 4622 41370
rect 4376 41316 4382 41318
rect 4438 41316 4462 41318
rect 4518 41316 4542 41318
rect 4598 41316 4622 41318
rect 4678 41316 4684 41318
rect 4376 41307 4684 41316
rect 7803 41372 8111 41381
rect 7803 41370 7809 41372
rect 7865 41370 7889 41372
rect 7945 41370 7969 41372
rect 8025 41370 8049 41372
rect 8105 41370 8111 41372
rect 7865 41318 7867 41370
rect 8047 41318 8049 41370
rect 7803 41316 7809 41318
rect 7865 41316 7889 41318
rect 7945 41316 7969 41318
rect 8025 41316 8049 41318
rect 8105 41316 8111 41318
rect 7803 41307 8111 41316
rect 11230 41372 11538 41381
rect 11230 41370 11236 41372
rect 11292 41370 11316 41372
rect 11372 41370 11396 41372
rect 11452 41370 11476 41372
rect 11532 41370 11538 41372
rect 11292 41318 11294 41370
rect 11474 41318 11476 41370
rect 11230 41316 11236 41318
rect 11292 41316 11316 41318
rect 11372 41316 11396 41318
rect 11452 41316 11476 41318
rect 11532 41316 11538 41318
rect 11230 41307 11538 41316
rect 14657 41372 14965 41381
rect 14657 41370 14663 41372
rect 14719 41370 14743 41372
rect 14799 41370 14823 41372
rect 14879 41370 14903 41372
rect 14959 41370 14965 41372
rect 14719 41318 14721 41370
rect 14901 41318 14903 41370
rect 14657 41316 14663 41318
rect 14719 41316 14743 41318
rect 14799 41316 14823 41318
rect 14879 41316 14903 41318
rect 14959 41316 14965 41318
rect 14657 41307 14965 41316
rect 2663 40828 2971 40837
rect 2663 40826 2669 40828
rect 2725 40826 2749 40828
rect 2805 40826 2829 40828
rect 2885 40826 2909 40828
rect 2965 40826 2971 40828
rect 2725 40774 2727 40826
rect 2907 40774 2909 40826
rect 2663 40772 2669 40774
rect 2725 40772 2749 40774
rect 2805 40772 2829 40774
rect 2885 40772 2909 40774
rect 2965 40772 2971 40774
rect 2663 40763 2971 40772
rect 6090 40828 6398 40837
rect 6090 40826 6096 40828
rect 6152 40826 6176 40828
rect 6232 40826 6256 40828
rect 6312 40826 6336 40828
rect 6392 40826 6398 40828
rect 6152 40774 6154 40826
rect 6334 40774 6336 40826
rect 6090 40772 6096 40774
rect 6152 40772 6176 40774
rect 6232 40772 6256 40774
rect 6312 40772 6336 40774
rect 6392 40772 6398 40774
rect 6090 40763 6398 40772
rect 9517 40828 9825 40837
rect 9517 40826 9523 40828
rect 9579 40826 9603 40828
rect 9659 40826 9683 40828
rect 9739 40826 9763 40828
rect 9819 40826 9825 40828
rect 9579 40774 9581 40826
rect 9761 40774 9763 40826
rect 9517 40772 9523 40774
rect 9579 40772 9603 40774
rect 9659 40772 9683 40774
rect 9739 40772 9763 40774
rect 9819 40772 9825 40774
rect 9517 40763 9825 40772
rect 12944 40828 13252 40837
rect 12944 40826 12950 40828
rect 13006 40826 13030 40828
rect 13086 40826 13110 40828
rect 13166 40826 13190 40828
rect 13246 40826 13252 40828
rect 13006 40774 13008 40826
rect 13188 40774 13190 40826
rect 12944 40772 12950 40774
rect 13006 40772 13030 40774
rect 13086 40772 13110 40774
rect 13166 40772 13190 40774
rect 13246 40772 13252 40774
rect 12944 40763 13252 40772
rect 4376 40284 4684 40293
rect 4376 40282 4382 40284
rect 4438 40282 4462 40284
rect 4518 40282 4542 40284
rect 4598 40282 4622 40284
rect 4678 40282 4684 40284
rect 4438 40230 4440 40282
rect 4620 40230 4622 40282
rect 4376 40228 4382 40230
rect 4438 40228 4462 40230
rect 4518 40228 4542 40230
rect 4598 40228 4622 40230
rect 4678 40228 4684 40230
rect 4376 40219 4684 40228
rect 7803 40284 8111 40293
rect 7803 40282 7809 40284
rect 7865 40282 7889 40284
rect 7945 40282 7969 40284
rect 8025 40282 8049 40284
rect 8105 40282 8111 40284
rect 7865 40230 7867 40282
rect 8047 40230 8049 40282
rect 7803 40228 7809 40230
rect 7865 40228 7889 40230
rect 7945 40228 7969 40230
rect 8025 40228 8049 40230
rect 8105 40228 8111 40230
rect 7803 40219 8111 40228
rect 11230 40284 11538 40293
rect 11230 40282 11236 40284
rect 11292 40282 11316 40284
rect 11372 40282 11396 40284
rect 11452 40282 11476 40284
rect 11532 40282 11538 40284
rect 11292 40230 11294 40282
rect 11474 40230 11476 40282
rect 11230 40228 11236 40230
rect 11292 40228 11316 40230
rect 11372 40228 11396 40230
rect 11452 40228 11476 40230
rect 11532 40228 11538 40230
rect 11230 40219 11538 40228
rect 14657 40284 14965 40293
rect 14657 40282 14663 40284
rect 14719 40282 14743 40284
rect 14799 40282 14823 40284
rect 14879 40282 14903 40284
rect 14959 40282 14965 40284
rect 14719 40230 14721 40282
rect 14901 40230 14903 40282
rect 14657 40228 14663 40230
rect 14719 40228 14743 40230
rect 14799 40228 14823 40230
rect 14879 40228 14903 40230
rect 14959 40228 14965 40230
rect 14657 40219 14965 40228
rect 2663 39740 2971 39749
rect 2663 39738 2669 39740
rect 2725 39738 2749 39740
rect 2805 39738 2829 39740
rect 2885 39738 2909 39740
rect 2965 39738 2971 39740
rect 2725 39686 2727 39738
rect 2907 39686 2909 39738
rect 2663 39684 2669 39686
rect 2725 39684 2749 39686
rect 2805 39684 2829 39686
rect 2885 39684 2909 39686
rect 2965 39684 2971 39686
rect 2663 39675 2971 39684
rect 6090 39740 6398 39749
rect 6090 39738 6096 39740
rect 6152 39738 6176 39740
rect 6232 39738 6256 39740
rect 6312 39738 6336 39740
rect 6392 39738 6398 39740
rect 6152 39686 6154 39738
rect 6334 39686 6336 39738
rect 6090 39684 6096 39686
rect 6152 39684 6176 39686
rect 6232 39684 6256 39686
rect 6312 39684 6336 39686
rect 6392 39684 6398 39686
rect 6090 39675 6398 39684
rect 9517 39740 9825 39749
rect 9517 39738 9523 39740
rect 9579 39738 9603 39740
rect 9659 39738 9683 39740
rect 9739 39738 9763 39740
rect 9819 39738 9825 39740
rect 9579 39686 9581 39738
rect 9761 39686 9763 39738
rect 9517 39684 9523 39686
rect 9579 39684 9603 39686
rect 9659 39684 9683 39686
rect 9739 39684 9763 39686
rect 9819 39684 9825 39686
rect 9517 39675 9825 39684
rect 12944 39740 13252 39749
rect 12944 39738 12950 39740
rect 13006 39738 13030 39740
rect 13086 39738 13110 39740
rect 13166 39738 13190 39740
rect 13246 39738 13252 39740
rect 13006 39686 13008 39738
rect 13188 39686 13190 39738
rect 12944 39684 12950 39686
rect 13006 39684 13030 39686
rect 13086 39684 13110 39686
rect 13166 39684 13190 39686
rect 13246 39684 13252 39686
rect 12944 39675 13252 39684
rect 4376 39196 4684 39205
rect 4376 39194 4382 39196
rect 4438 39194 4462 39196
rect 4518 39194 4542 39196
rect 4598 39194 4622 39196
rect 4678 39194 4684 39196
rect 4438 39142 4440 39194
rect 4620 39142 4622 39194
rect 4376 39140 4382 39142
rect 4438 39140 4462 39142
rect 4518 39140 4542 39142
rect 4598 39140 4622 39142
rect 4678 39140 4684 39142
rect 4376 39131 4684 39140
rect 7803 39196 8111 39205
rect 7803 39194 7809 39196
rect 7865 39194 7889 39196
rect 7945 39194 7969 39196
rect 8025 39194 8049 39196
rect 8105 39194 8111 39196
rect 7865 39142 7867 39194
rect 8047 39142 8049 39194
rect 7803 39140 7809 39142
rect 7865 39140 7889 39142
rect 7945 39140 7969 39142
rect 8025 39140 8049 39142
rect 8105 39140 8111 39142
rect 7803 39131 8111 39140
rect 11230 39196 11538 39205
rect 11230 39194 11236 39196
rect 11292 39194 11316 39196
rect 11372 39194 11396 39196
rect 11452 39194 11476 39196
rect 11532 39194 11538 39196
rect 11292 39142 11294 39194
rect 11474 39142 11476 39194
rect 11230 39140 11236 39142
rect 11292 39140 11316 39142
rect 11372 39140 11396 39142
rect 11452 39140 11476 39142
rect 11532 39140 11538 39142
rect 11230 39131 11538 39140
rect 14657 39196 14965 39205
rect 14657 39194 14663 39196
rect 14719 39194 14743 39196
rect 14799 39194 14823 39196
rect 14879 39194 14903 39196
rect 14959 39194 14965 39196
rect 14719 39142 14721 39194
rect 14901 39142 14903 39194
rect 14657 39140 14663 39142
rect 14719 39140 14743 39142
rect 14799 39140 14823 39142
rect 14879 39140 14903 39142
rect 14959 39140 14965 39142
rect 14657 39131 14965 39140
rect 2663 38652 2971 38661
rect 2663 38650 2669 38652
rect 2725 38650 2749 38652
rect 2805 38650 2829 38652
rect 2885 38650 2909 38652
rect 2965 38650 2971 38652
rect 2725 38598 2727 38650
rect 2907 38598 2909 38650
rect 2663 38596 2669 38598
rect 2725 38596 2749 38598
rect 2805 38596 2829 38598
rect 2885 38596 2909 38598
rect 2965 38596 2971 38598
rect 2663 38587 2971 38596
rect 6090 38652 6398 38661
rect 6090 38650 6096 38652
rect 6152 38650 6176 38652
rect 6232 38650 6256 38652
rect 6312 38650 6336 38652
rect 6392 38650 6398 38652
rect 6152 38598 6154 38650
rect 6334 38598 6336 38650
rect 6090 38596 6096 38598
rect 6152 38596 6176 38598
rect 6232 38596 6256 38598
rect 6312 38596 6336 38598
rect 6392 38596 6398 38598
rect 6090 38587 6398 38596
rect 9517 38652 9825 38661
rect 9517 38650 9523 38652
rect 9579 38650 9603 38652
rect 9659 38650 9683 38652
rect 9739 38650 9763 38652
rect 9819 38650 9825 38652
rect 9579 38598 9581 38650
rect 9761 38598 9763 38650
rect 9517 38596 9523 38598
rect 9579 38596 9603 38598
rect 9659 38596 9683 38598
rect 9739 38596 9763 38598
rect 9819 38596 9825 38598
rect 9517 38587 9825 38596
rect 12944 38652 13252 38661
rect 12944 38650 12950 38652
rect 13006 38650 13030 38652
rect 13086 38650 13110 38652
rect 13166 38650 13190 38652
rect 13246 38650 13252 38652
rect 13006 38598 13008 38650
rect 13188 38598 13190 38650
rect 12944 38596 12950 38598
rect 13006 38596 13030 38598
rect 13086 38596 13110 38598
rect 13166 38596 13190 38598
rect 13246 38596 13252 38598
rect 12944 38587 13252 38596
rect 4376 38108 4684 38117
rect 4376 38106 4382 38108
rect 4438 38106 4462 38108
rect 4518 38106 4542 38108
rect 4598 38106 4622 38108
rect 4678 38106 4684 38108
rect 4438 38054 4440 38106
rect 4620 38054 4622 38106
rect 4376 38052 4382 38054
rect 4438 38052 4462 38054
rect 4518 38052 4542 38054
rect 4598 38052 4622 38054
rect 4678 38052 4684 38054
rect 4376 38043 4684 38052
rect 7803 38108 8111 38117
rect 7803 38106 7809 38108
rect 7865 38106 7889 38108
rect 7945 38106 7969 38108
rect 8025 38106 8049 38108
rect 8105 38106 8111 38108
rect 7865 38054 7867 38106
rect 8047 38054 8049 38106
rect 7803 38052 7809 38054
rect 7865 38052 7889 38054
rect 7945 38052 7969 38054
rect 8025 38052 8049 38054
rect 8105 38052 8111 38054
rect 7803 38043 8111 38052
rect 11230 38108 11538 38117
rect 11230 38106 11236 38108
rect 11292 38106 11316 38108
rect 11372 38106 11396 38108
rect 11452 38106 11476 38108
rect 11532 38106 11538 38108
rect 11292 38054 11294 38106
rect 11474 38054 11476 38106
rect 11230 38052 11236 38054
rect 11292 38052 11316 38054
rect 11372 38052 11396 38054
rect 11452 38052 11476 38054
rect 11532 38052 11538 38054
rect 11230 38043 11538 38052
rect 14657 38108 14965 38117
rect 14657 38106 14663 38108
rect 14719 38106 14743 38108
rect 14799 38106 14823 38108
rect 14879 38106 14903 38108
rect 14959 38106 14965 38108
rect 14719 38054 14721 38106
rect 14901 38054 14903 38106
rect 14657 38052 14663 38054
rect 14719 38052 14743 38054
rect 14799 38052 14823 38054
rect 14879 38052 14903 38054
rect 14959 38052 14965 38054
rect 14657 38043 14965 38052
rect 2663 37564 2971 37573
rect 2663 37562 2669 37564
rect 2725 37562 2749 37564
rect 2805 37562 2829 37564
rect 2885 37562 2909 37564
rect 2965 37562 2971 37564
rect 2725 37510 2727 37562
rect 2907 37510 2909 37562
rect 2663 37508 2669 37510
rect 2725 37508 2749 37510
rect 2805 37508 2829 37510
rect 2885 37508 2909 37510
rect 2965 37508 2971 37510
rect 2663 37499 2971 37508
rect 6090 37564 6398 37573
rect 6090 37562 6096 37564
rect 6152 37562 6176 37564
rect 6232 37562 6256 37564
rect 6312 37562 6336 37564
rect 6392 37562 6398 37564
rect 6152 37510 6154 37562
rect 6334 37510 6336 37562
rect 6090 37508 6096 37510
rect 6152 37508 6176 37510
rect 6232 37508 6256 37510
rect 6312 37508 6336 37510
rect 6392 37508 6398 37510
rect 6090 37499 6398 37508
rect 9517 37564 9825 37573
rect 9517 37562 9523 37564
rect 9579 37562 9603 37564
rect 9659 37562 9683 37564
rect 9739 37562 9763 37564
rect 9819 37562 9825 37564
rect 9579 37510 9581 37562
rect 9761 37510 9763 37562
rect 9517 37508 9523 37510
rect 9579 37508 9603 37510
rect 9659 37508 9683 37510
rect 9739 37508 9763 37510
rect 9819 37508 9825 37510
rect 9517 37499 9825 37508
rect 12944 37564 13252 37573
rect 12944 37562 12950 37564
rect 13006 37562 13030 37564
rect 13086 37562 13110 37564
rect 13166 37562 13190 37564
rect 13246 37562 13252 37564
rect 13006 37510 13008 37562
rect 13188 37510 13190 37562
rect 12944 37508 12950 37510
rect 13006 37508 13030 37510
rect 13086 37508 13110 37510
rect 13166 37508 13190 37510
rect 13246 37508 13252 37510
rect 12944 37499 13252 37508
rect 4376 37020 4684 37029
rect 4376 37018 4382 37020
rect 4438 37018 4462 37020
rect 4518 37018 4542 37020
rect 4598 37018 4622 37020
rect 4678 37018 4684 37020
rect 4438 36966 4440 37018
rect 4620 36966 4622 37018
rect 4376 36964 4382 36966
rect 4438 36964 4462 36966
rect 4518 36964 4542 36966
rect 4598 36964 4622 36966
rect 4678 36964 4684 36966
rect 4376 36955 4684 36964
rect 7803 37020 8111 37029
rect 7803 37018 7809 37020
rect 7865 37018 7889 37020
rect 7945 37018 7969 37020
rect 8025 37018 8049 37020
rect 8105 37018 8111 37020
rect 7865 36966 7867 37018
rect 8047 36966 8049 37018
rect 7803 36964 7809 36966
rect 7865 36964 7889 36966
rect 7945 36964 7969 36966
rect 8025 36964 8049 36966
rect 8105 36964 8111 36966
rect 7803 36955 8111 36964
rect 11230 37020 11538 37029
rect 11230 37018 11236 37020
rect 11292 37018 11316 37020
rect 11372 37018 11396 37020
rect 11452 37018 11476 37020
rect 11532 37018 11538 37020
rect 11292 36966 11294 37018
rect 11474 36966 11476 37018
rect 11230 36964 11236 36966
rect 11292 36964 11316 36966
rect 11372 36964 11396 36966
rect 11452 36964 11476 36966
rect 11532 36964 11538 36966
rect 11230 36955 11538 36964
rect 14657 37020 14965 37029
rect 14657 37018 14663 37020
rect 14719 37018 14743 37020
rect 14799 37018 14823 37020
rect 14879 37018 14903 37020
rect 14959 37018 14965 37020
rect 14719 36966 14721 37018
rect 14901 36966 14903 37018
rect 14657 36964 14663 36966
rect 14719 36964 14743 36966
rect 14799 36964 14823 36966
rect 14879 36964 14903 36966
rect 14959 36964 14965 36966
rect 14657 36955 14965 36964
rect 2663 36476 2971 36485
rect 2663 36474 2669 36476
rect 2725 36474 2749 36476
rect 2805 36474 2829 36476
rect 2885 36474 2909 36476
rect 2965 36474 2971 36476
rect 2725 36422 2727 36474
rect 2907 36422 2909 36474
rect 2663 36420 2669 36422
rect 2725 36420 2749 36422
rect 2805 36420 2829 36422
rect 2885 36420 2909 36422
rect 2965 36420 2971 36422
rect 2663 36411 2971 36420
rect 6090 36476 6398 36485
rect 6090 36474 6096 36476
rect 6152 36474 6176 36476
rect 6232 36474 6256 36476
rect 6312 36474 6336 36476
rect 6392 36474 6398 36476
rect 6152 36422 6154 36474
rect 6334 36422 6336 36474
rect 6090 36420 6096 36422
rect 6152 36420 6176 36422
rect 6232 36420 6256 36422
rect 6312 36420 6336 36422
rect 6392 36420 6398 36422
rect 6090 36411 6398 36420
rect 9517 36476 9825 36485
rect 9517 36474 9523 36476
rect 9579 36474 9603 36476
rect 9659 36474 9683 36476
rect 9739 36474 9763 36476
rect 9819 36474 9825 36476
rect 9579 36422 9581 36474
rect 9761 36422 9763 36474
rect 9517 36420 9523 36422
rect 9579 36420 9603 36422
rect 9659 36420 9683 36422
rect 9739 36420 9763 36422
rect 9819 36420 9825 36422
rect 9517 36411 9825 36420
rect 12944 36476 13252 36485
rect 12944 36474 12950 36476
rect 13006 36474 13030 36476
rect 13086 36474 13110 36476
rect 13166 36474 13190 36476
rect 13246 36474 13252 36476
rect 13006 36422 13008 36474
rect 13188 36422 13190 36474
rect 12944 36420 12950 36422
rect 13006 36420 13030 36422
rect 13086 36420 13110 36422
rect 13166 36420 13190 36422
rect 13246 36420 13252 36422
rect 12944 36411 13252 36420
rect 14464 36032 14516 36038
rect 14464 35974 14516 35980
rect 4376 35932 4684 35941
rect 4376 35930 4382 35932
rect 4438 35930 4462 35932
rect 4518 35930 4542 35932
rect 4598 35930 4622 35932
rect 4678 35930 4684 35932
rect 4438 35878 4440 35930
rect 4620 35878 4622 35930
rect 4376 35876 4382 35878
rect 4438 35876 4462 35878
rect 4518 35876 4542 35878
rect 4598 35876 4622 35878
rect 4678 35876 4684 35878
rect 4376 35867 4684 35876
rect 7803 35932 8111 35941
rect 7803 35930 7809 35932
rect 7865 35930 7889 35932
rect 7945 35930 7969 35932
rect 8025 35930 8049 35932
rect 8105 35930 8111 35932
rect 7865 35878 7867 35930
rect 8047 35878 8049 35930
rect 7803 35876 7809 35878
rect 7865 35876 7889 35878
rect 7945 35876 7969 35878
rect 8025 35876 8049 35878
rect 8105 35876 8111 35878
rect 7803 35867 8111 35876
rect 11230 35932 11538 35941
rect 11230 35930 11236 35932
rect 11292 35930 11316 35932
rect 11372 35930 11396 35932
rect 11452 35930 11476 35932
rect 11532 35930 11538 35932
rect 11292 35878 11294 35930
rect 11474 35878 11476 35930
rect 11230 35876 11236 35878
rect 11292 35876 11316 35878
rect 11372 35876 11396 35878
rect 11452 35876 11476 35878
rect 11532 35876 11538 35878
rect 11230 35867 11538 35876
rect 14476 35737 14504 35974
rect 14657 35932 14965 35941
rect 14657 35930 14663 35932
rect 14719 35930 14743 35932
rect 14799 35930 14823 35932
rect 14879 35930 14903 35932
rect 14959 35930 14965 35932
rect 14719 35878 14721 35930
rect 14901 35878 14903 35930
rect 14657 35876 14663 35878
rect 14719 35876 14743 35878
rect 14799 35876 14823 35878
rect 14879 35876 14903 35878
rect 14959 35876 14965 35878
rect 14657 35867 14965 35876
rect 14462 35728 14518 35737
rect 14462 35663 14518 35672
rect 2663 35388 2971 35397
rect 2663 35386 2669 35388
rect 2725 35386 2749 35388
rect 2805 35386 2829 35388
rect 2885 35386 2909 35388
rect 2965 35386 2971 35388
rect 2725 35334 2727 35386
rect 2907 35334 2909 35386
rect 2663 35332 2669 35334
rect 2725 35332 2749 35334
rect 2805 35332 2829 35334
rect 2885 35332 2909 35334
rect 2965 35332 2971 35334
rect 2663 35323 2971 35332
rect 6090 35388 6398 35397
rect 6090 35386 6096 35388
rect 6152 35386 6176 35388
rect 6232 35386 6256 35388
rect 6312 35386 6336 35388
rect 6392 35386 6398 35388
rect 6152 35334 6154 35386
rect 6334 35334 6336 35386
rect 6090 35332 6096 35334
rect 6152 35332 6176 35334
rect 6232 35332 6256 35334
rect 6312 35332 6336 35334
rect 6392 35332 6398 35334
rect 6090 35323 6398 35332
rect 9517 35388 9825 35397
rect 9517 35386 9523 35388
rect 9579 35386 9603 35388
rect 9659 35386 9683 35388
rect 9739 35386 9763 35388
rect 9819 35386 9825 35388
rect 9579 35334 9581 35386
rect 9761 35334 9763 35386
rect 9517 35332 9523 35334
rect 9579 35332 9603 35334
rect 9659 35332 9683 35334
rect 9739 35332 9763 35334
rect 9819 35332 9825 35334
rect 9517 35323 9825 35332
rect 12944 35388 13252 35397
rect 12944 35386 12950 35388
rect 13006 35386 13030 35388
rect 13086 35386 13110 35388
rect 13166 35386 13190 35388
rect 13246 35386 13252 35388
rect 13006 35334 13008 35386
rect 13188 35334 13190 35386
rect 12944 35332 12950 35334
rect 13006 35332 13030 35334
rect 13086 35332 13110 35334
rect 13166 35332 13190 35334
rect 13246 35332 13252 35334
rect 12944 35323 13252 35332
rect 4376 34844 4684 34853
rect 4376 34842 4382 34844
rect 4438 34842 4462 34844
rect 4518 34842 4542 34844
rect 4598 34842 4622 34844
rect 4678 34842 4684 34844
rect 4438 34790 4440 34842
rect 4620 34790 4622 34842
rect 4376 34788 4382 34790
rect 4438 34788 4462 34790
rect 4518 34788 4542 34790
rect 4598 34788 4622 34790
rect 4678 34788 4684 34790
rect 4376 34779 4684 34788
rect 7803 34844 8111 34853
rect 7803 34842 7809 34844
rect 7865 34842 7889 34844
rect 7945 34842 7969 34844
rect 8025 34842 8049 34844
rect 8105 34842 8111 34844
rect 7865 34790 7867 34842
rect 8047 34790 8049 34842
rect 7803 34788 7809 34790
rect 7865 34788 7889 34790
rect 7945 34788 7969 34790
rect 8025 34788 8049 34790
rect 8105 34788 8111 34790
rect 7803 34779 8111 34788
rect 11230 34844 11538 34853
rect 11230 34842 11236 34844
rect 11292 34842 11316 34844
rect 11372 34842 11396 34844
rect 11452 34842 11476 34844
rect 11532 34842 11538 34844
rect 11292 34790 11294 34842
rect 11474 34790 11476 34842
rect 11230 34788 11236 34790
rect 11292 34788 11316 34790
rect 11372 34788 11396 34790
rect 11452 34788 11476 34790
rect 11532 34788 11538 34790
rect 11230 34779 11538 34788
rect 14657 34844 14965 34853
rect 14657 34842 14663 34844
rect 14719 34842 14743 34844
rect 14799 34842 14823 34844
rect 14879 34842 14903 34844
rect 14959 34842 14965 34844
rect 14719 34790 14721 34842
rect 14901 34790 14903 34842
rect 14657 34788 14663 34790
rect 14719 34788 14743 34790
rect 14799 34788 14823 34790
rect 14879 34788 14903 34790
rect 14959 34788 14965 34790
rect 14657 34779 14965 34788
rect 2663 34300 2971 34309
rect 2663 34298 2669 34300
rect 2725 34298 2749 34300
rect 2805 34298 2829 34300
rect 2885 34298 2909 34300
rect 2965 34298 2971 34300
rect 2725 34246 2727 34298
rect 2907 34246 2909 34298
rect 2663 34244 2669 34246
rect 2725 34244 2749 34246
rect 2805 34244 2829 34246
rect 2885 34244 2909 34246
rect 2965 34244 2971 34246
rect 2663 34235 2971 34244
rect 6090 34300 6398 34309
rect 6090 34298 6096 34300
rect 6152 34298 6176 34300
rect 6232 34298 6256 34300
rect 6312 34298 6336 34300
rect 6392 34298 6398 34300
rect 6152 34246 6154 34298
rect 6334 34246 6336 34298
rect 6090 34244 6096 34246
rect 6152 34244 6176 34246
rect 6232 34244 6256 34246
rect 6312 34244 6336 34246
rect 6392 34244 6398 34246
rect 6090 34235 6398 34244
rect 9517 34300 9825 34309
rect 9517 34298 9523 34300
rect 9579 34298 9603 34300
rect 9659 34298 9683 34300
rect 9739 34298 9763 34300
rect 9819 34298 9825 34300
rect 9579 34246 9581 34298
rect 9761 34246 9763 34298
rect 9517 34244 9523 34246
rect 9579 34244 9603 34246
rect 9659 34244 9683 34246
rect 9739 34244 9763 34246
rect 9819 34244 9825 34246
rect 9517 34235 9825 34244
rect 12944 34300 13252 34309
rect 12944 34298 12950 34300
rect 13006 34298 13030 34300
rect 13086 34298 13110 34300
rect 13166 34298 13190 34300
rect 13246 34298 13252 34300
rect 13006 34246 13008 34298
rect 13188 34246 13190 34298
rect 12944 34244 12950 34246
rect 13006 34244 13030 34246
rect 13086 34244 13110 34246
rect 13166 34244 13190 34246
rect 13246 34244 13252 34246
rect 12944 34235 13252 34244
rect 4376 33756 4684 33765
rect 4376 33754 4382 33756
rect 4438 33754 4462 33756
rect 4518 33754 4542 33756
rect 4598 33754 4622 33756
rect 4678 33754 4684 33756
rect 4438 33702 4440 33754
rect 4620 33702 4622 33754
rect 4376 33700 4382 33702
rect 4438 33700 4462 33702
rect 4518 33700 4542 33702
rect 4598 33700 4622 33702
rect 4678 33700 4684 33702
rect 4376 33691 4684 33700
rect 7803 33756 8111 33765
rect 7803 33754 7809 33756
rect 7865 33754 7889 33756
rect 7945 33754 7969 33756
rect 8025 33754 8049 33756
rect 8105 33754 8111 33756
rect 7865 33702 7867 33754
rect 8047 33702 8049 33754
rect 7803 33700 7809 33702
rect 7865 33700 7889 33702
rect 7945 33700 7969 33702
rect 8025 33700 8049 33702
rect 8105 33700 8111 33702
rect 7803 33691 8111 33700
rect 11230 33756 11538 33765
rect 11230 33754 11236 33756
rect 11292 33754 11316 33756
rect 11372 33754 11396 33756
rect 11452 33754 11476 33756
rect 11532 33754 11538 33756
rect 11292 33702 11294 33754
rect 11474 33702 11476 33754
rect 11230 33700 11236 33702
rect 11292 33700 11316 33702
rect 11372 33700 11396 33702
rect 11452 33700 11476 33702
rect 11532 33700 11538 33702
rect 11230 33691 11538 33700
rect 14657 33756 14965 33765
rect 14657 33754 14663 33756
rect 14719 33754 14743 33756
rect 14799 33754 14823 33756
rect 14879 33754 14903 33756
rect 14959 33754 14965 33756
rect 14719 33702 14721 33754
rect 14901 33702 14903 33754
rect 14657 33700 14663 33702
rect 14719 33700 14743 33702
rect 14799 33700 14823 33702
rect 14879 33700 14903 33702
rect 14959 33700 14965 33702
rect 14657 33691 14965 33700
rect 2663 33212 2971 33221
rect 2663 33210 2669 33212
rect 2725 33210 2749 33212
rect 2805 33210 2829 33212
rect 2885 33210 2909 33212
rect 2965 33210 2971 33212
rect 2725 33158 2727 33210
rect 2907 33158 2909 33210
rect 2663 33156 2669 33158
rect 2725 33156 2749 33158
rect 2805 33156 2829 33158
rect 2885 33156 2909 33158
rect 2965 33156 2971 33158
rect 2663 33147 2971 33156
rect 6090 33212 6398 33221
rect 6090 33210 6096 33212
rect 6152 33210 6176 33212
rect 6232 33210 6256 33212
rect 6312 33210 6336 33212
rect 6392 33210 6398 33212
rect 6152 33158 6154 33210
rect 6334 33158 6336 33210
rect 6090 33156 6096 33158
rect 6152 33156 6176 33158
rect 6232 33156 6256 33158
rect 6312 33156 6336 33158
rect 6392 33156 6398 33158
rect 6090 33147 6398 33156
rect 9517 33212 9825 33221
rect 9517 33210 9523 33212
rect 9579 33210 9603 33212
rect 9659 33210 9683 33212
rect 9739 33210 9763 33212
rect 9819 33210 9825 33212
rect 9579 33158 9581 33210
rect 9761 33158 9763 33210
rect 9517 33156 9523 33158
rect 9579 33156 9603 33158
rect 9659 33156 9683 33158
rect 9739 33156 9763 33158
rect 9819 33156 9825 33158
rect 9517 33147 9825 33156
rect 12944 33212 13252 33221
rect 12944 33210 12950 33212
rect 13006 33210 13030 33212
rect 13086 33210 13110 33212
rect 13166 33210 13190 33212
rect 13246 33210 13252 33212
rect 13006 33158 13008 33210
rect 13188 33158 13190 33210
rect 12944 33156 12950 33158
rect 13006 33156 13030 33158
rect 13086 33156 13110 33158
rect 13166 33156 13190 33158
rect 13246 33156 13252 33158
rect 12944 33147 13252 33156
rect 4376 32668 4684 32677
rect 4376 32666 4382 32668
rect 4438 32666 4462 32668
rect 4518 32666 4542 32668
rect 4598 32666 4622 32668
rect 4678 32666 4684 32668
rect 4438 32614 4440 32666
rect 4620 32614 4622 32666
rect 4376 32612 4382 32614
rect 4438 32612 4462 32614
rect 4518 32612 4542 32614
rect 4598 32612 4622 32614
rect 4678 32612 4684 32614
rect 4376 32603 4684 32612
rect 7803 32668 8111 32677
rect 7803 32666 7809 32668
rect 7865 32666 7889 32668
rect 7945 32666 7969 32668
rect 8025 32666 8049 32668
rect 8105 32666 8111 32668
rect 7865 32614 7867 32666
rect 8047 32614 8049 32666
rect 7803 32612 7809 32614
rect 7865 32612 7889 32614
rect 7945 32612 7969 32614
rect 8025 32612 8049 32614
rect 8105 32612 8111 32614
rect 7803 32603 8111 32612
rect 11230 32668 11538 32677
rect 11230 32666 11236 32668
rect 11292 32666 11316 32668
rect 11372 32666 11396 32668
rect 11452 32666 11476 32668
rect 11532 32666 11538 32668
rect 11292 32614 11294 32666
rect 11474 32614 11476 32666
rect 11230 32612 11236 32614
rect 11292 32612 11316 32614
rect 11372 32612 11396 32614
rect 11452 32612 11476 32614
rect 11532 32612 11538 32614
rect 11230 32603 11538 32612
rect 14657 32668 14965 32677
rect 14657 32666 14663 32668
rect 14719 32666 14743 32668
rect 14799 32666 14823 32668
rect 14879 32666 14903 32668
rect 14959 32666 14965 32668
rect 14719 32614 14721 32666
rect 14901 32614 14903 32666
rect 14657 32612 14663 32614
rect 14719 32612 14743 32614
rect 14799 32612 14823 32614
rect 14879 32612 14903 32614
rect 14959 32612 14965 32614
rect 14657 32603 14965 32612
rect 2663 32124 2971 32133
rect 2663 32122 2669 32124
rect 2725 32122 2749 32124
rect 2805 32122 2829 32124
rect 2885 32122 2909 32124
rect 2965 32122 2971 32124
rect 2725 32070 2727 32122
rect 2907 32070 2909 32122
rect 2663 32068 2669 32070
rect 2725 32068 2749 32070
rect 2805 32068 2829 32070
rect 2885 32068 2909 32070
rect 2965 32068 2971 32070
rect 2663 32059 2971 32068
rect 6090 32124 6398 32133
rect 6090 32122 6096 32124
rect 6152 32122 6176 32124
rect 6232 32122 6256 32124
rect 6312 32122 6336 32124
rect 6392 32122 6398 32124
rect 6152 32070 6154 32122
rect 6334 32070 6336 32122
rect 6090 32068 6096 32070
rect 6152 32068 6176 32070
rect 6232 32068 6256 32070
rect 6312 32068 6336 32070
rect 6392 32068 6398 32070
rect 6090 32059 6398 32068
rect 9517 32124 9825 32133
rect 9517 32122 9523 32124
rect 9579 32122 9603 32124
rect 9659 32122 9683 32124
rect 9739 32122 9763 32124
rect 9819 32122 9825 32124
rect 9579 32070 9581 32122
rect 9761 32070 9763 32122
rect 9517 32068 9523 32070
rect 9579 32068 9603 32070
rect 9659 32068 9683 32070
rect 9739 32068 9763 32070
rect 9819 32068 9825 32070
rect 9517 32059 9825 32068
rect 12944 32124 13252 32133
rect 12944 32122 12950 32124
rect 13006 32122 13030 32124
rect 13086 32122 13110 32124
rect 13166 32122 13190 32124
rect 13246 32122 13252 32124
rect 13006 32070 13008 32122
rect 13188 32070 13190 32122
rect 12944 32068 12950 32070
rect 13006 32068 13030 32070
rect 13086 32068 13110 32070
rect 13166 32068 13190 32070
rect 13246 32068 13252 32070
rect 12944 32059 13252 32068
rect 4376 31580 4684 31589
rect 4376 31578 4382 31580
rect 4438 31578 4462 31580
rect 4518 31578 4542 31580
rect 4598 31578 4622 31580
rect 4678 31578 4684 31580
rect 4438 31526 4440 31578
rect 4620 31526 4622 31578
rect 4376 31524 4382 31526
rect 4438 31524 4462 31526
rect 4518 31524 4542 31526
rect 4598 31524 4622 31526
rect 4678 31524 4684 31526
rect 4376 31515 4684 31524
rect 7803 31580 8111 31589
rect 7803 31578 7809 31580
rect 7865 31578 7889 31580
rect 7945 31578 7969 31580
rect 8025 31578 8049 31580
rect 8105 31578 8111 31580
rect 7865 31526 7867 31578
rect 8047 31526 8049 31578
rect 7803 31524 7809 31526
rect 7865 31524 7889 31526
rect 7945 31524 7969 31526
rect 8025 31524 8049 31526
rect 8105 31524 8111 31526
rect 7803 31515 8111 31524
rect 11230 31580 11538 31589
rect 11230 31578 11236 31580
rect 11292 31578 11316 31580
rect 11372 31578 11396 31580
rect 11452 31578 11476 31580
rect 11532 31578 11538 31580
rect 11292 31526 11294 31578
rect 11474 31526 11476 31578
rect 11230 31524 11236 31526
rect 11292 31524 11316 31526
rect 11372 31524 11396 31526
rect 11452 31524 11476 31526
rect 11532 31524 11538 31526
rect 11230 31515 11538 31524
rect 14657 31580 14965 31589
rect 14657 31578 14663 31580
rect 14719 31578 14743 31580
rect 14799 31578 14823 31580
rect 14879 31578 14903 31580
rect 14959 31578 14965 31580
rect 14719 31526 14721 31578
rect 14901 31526 14903 31578
rect 14657 31524 14663 31526
rect 14719 31524 14743 31526
rect 14799 31524 14823 31526
rect 14879 31524 14903 31526
rect 14959 31524 14965 31526
rect 14657 31515 14965 31524
rect 2663 31036 2971 31045
rect 2663 31034 2669 31036
rect 2725 31034 2749 31036
rect 2805 31034 2829 31036
rect 2885 31034 2909 31036
rect 2965 31034 2971 31036
rect 2725 30982 2727 31034
rect 2907 30982 2909 31034
rect 2663 30980 2669 30982
rect 2725 30980 2749 30982
rect 2805 30980 2829 30982
rect 2885 30980 2909 30982
rect 2965 30980 2971 30982
rect 2663 30971 2971 30980
rect 6090 31036 6398 31045
rect 6090 31034 6096 31036
rect 6152 31034 6176 31036
rect 6232 31034 6256 31036
rect 6312 31034 6336 31036
rect 6392 31034 6398 31036
rect 6152 30982 6154 31034
rect 6334 30982 6336 31034
rect 6090 30980 6096 30982
rect 6152 30980 6176 30982
rect 6232 30980 6256 30982
rect 6312 30980 6336 30982
rect 6392 30980 6398 30982
rect 6090 30971 6398 30980
rect 9517 31036 9825 31045
rect 9517 31034 9523 31036
rect 9579 31034 9603 31036
rect 9659 31034 9683 31036
rect 9739 31034 9763 31036
rect 9819 31034 9825 31036
rect 9579 30982 9581 31034
rect 9761 30982 9763 31034
rect 9517 30980 9523 30982
rect 9579 30980 9603 30982
rect 9659 30980 9683 30982
rect 9739 30980 9763 30982
rect 9819 30980 9825 30982
rect 9517 30971 9825 30980
rect 12944 31036 13252 31045
rect 12944 31034 12950 31036
rect 13006 31034 13030 31036
rect 13086 31034 13110 31036
rect 13166 31034 13190 31036
rect 13246 31034 13252 31036
rect 13006 30982 13008 31034
rect 13188 30982 13190 31034
rect 12944 30980 12950 30982
rect 13006 30980 13030 30982
rect 13086 30980 13110 30982
rect 13166 30980 13190 30982
rect 13246 30980 13252 30982
rect 12944 30971 13252 30980
rect 4376 30492 4684 30501
rect 4376 30490 4382 30492
rect 4438 30490 4462 30492
rect 4518 30490 4542 30492
rect 4598 30490 4622 30492
rect 4678 30490 4684 30492
rect 4438 30438 4440 30490
rect 4620 30438 4622 30490
rect 4376 30436 4382 30438
rect 4438 30436 4462 30438
rect 4518 30436 4542 30438
rect 4598 30436 4622 30438
rect 4678 30436 4684 30438
rect 4376 30427 4684 30436
rect 7803 30492 8111 30501
rect 7803 30490 7809 30492
rect 7865 30490 7889 30492
rect 7945 30490 7969 30492
rect 8025 30490 8049 30492
rect 8105 30490 8111 30492
rect 7865 30438 7867 30490
rect 8047 30438 8049 30490
rect 7803 30436 7809 30438
rect 7865 30436 7889 30438
rect 7945 30436 7969 30438
rect 8025 30436 8049 30438
rect 8105 30436 8111 30438
rect 7803 30427 8111 30436
rect 11230 30492 11538 30501
rect 11230 30490 11236 30492
rect 11292 30490 11316 30492
rect 11372 30490 11396 30492
rect 11452 30490 11476 30492
rect 11532 30490 11538 30492
rect 11292 30438 11294 30490
rect 11474 30438 11476 30490
rect 11230 30436 11236 30438
rect 11292 30436 11316 30438
rect 11372 30436 11396 30438
rect 11452 30436 11476 30438
rect 11532 30436 11538 30438
rect 11230 30427 11538 30436
rect 14657 30492 14965 30501
rect 14657 30490 14663 30492
rect 14719 30490 14743 30492
rect 14799 30490 14823 30492
rect 14879 30490 14903 30492
rect 14959 30490 14965 30492
rect 14719 30438 14721 30490
rect 14901 30438 14903 30490
rect 14657 30436 14663 30438
rect 14719 30436 14743 30438
rect 14799 30436 14823 30438
rect 14879 30436 14903 30438
rect 14959 30436 14965 30438
rect 14657 30427 14965 30436
rect 2663 29948 2971 29957
rect 2663 29946 2669 29948
rect 2725 29946 2749 29948
rect 2805 29946 2829 29948
rect 2885 29946 2909 29948
rect 2965 29946 2971 29948
rect 2725 29894 2727 29946
rect 2907 29894 2909 29946
rect 2663 29892 2669 29894
rect 2725 29892 2749 29894
rect 2805 29892 2829 29894
rect 2885 29892 2909 29894
rect 2965 29892 2971 29894
rect 2663 29883 2971 29892
rect 6090 29948 6398 29957
rect 6090 29946 6096 29948
rect 6152 29946 6176 29948
rect 6232 29946 6256 29948
rect 6312 29946 6336 29948
rect 6392 29946 6398 29948
rect 6152 29894 6154 29946
rect 6334 29894 6336 29946
rect 6090 29892 6096 29894
rect 6152 29892 6176 29894
rect 6232 29892 6256 29894
rect 6312 29892 6336 29894
rect 6392 29892 6398 29894
rect 6090 29883 6398 29892
rect 9517 29948 9825 29957
rect 9517 29946 9523 29948
rect 9579 29946 9603 29948
rect 9659 29946 9683 29948
rect 9739 29946 9763 29948
rect 9819 29946 9825 29948
rect 9579 29894 9581 29946
rect 9761 29894 9763 29946
rect 9517 29892 9523 29894
rect 9579 29892 9603 29894
rect 9659 29892 9683 29894
rect 9739 29892 9763 29894
rect 9819 29892 9825 29894
rect 9517 29883 9825 29892
rect 12944 29948 13252 29957
rect 12944 29946 12950 29948
rect 13006 29946 13030 29948
rect 13086 29946 13110 29948
rect 13166 29946 13190 29948
rect 13246 29946 13252 29948
rect 13006 29894 13008 29946
rect 13188 29894 13190 29946
rect 12944 29892 12950 29894
rect 13006 29892 13030 29894
rect 13086 29892 13110 29894
rect 13166 29892 13190 29894
rect 13246 29892 13252 29894
rect 12944 29883 13252 29892
rect 4376 29404 4684 29413
rect 4376 29402 4382 29404
rect 4438 29402 4462 29404
rect 4518 29402 4542 29404
rect 4598 29402 4622 29404
rect 4678 29402 4684 29404
rect 4438 29350 4440 29402
rect 4620 29350 4622 29402
rect 4376 29348 4382 29350
rect 4438 29348 4462 29350
rect 4518 29348 4542 29350
rect 4598 29348 4622 29350
rect 4678 29348 4684 29350
rect 4376 29339 4684 29348
rect 7803 29404 8111 29413
rect 7803 29402 7809 29404
rect 7865 29402 7889 29404
rect 7945 29402 7969 29404
rect 8025 29402 8049 29404
rect 8105 29402 8111 29404
rect 7865 29350 7867 29402
rect 8047 29350 8049 29402
rect 7803 29348 7809 29350
rect 7865 29348 7889 29350
rect 7945 29348 7969 29350
rect 8025 29348 8049 29350
rect 8105 29348 8111 29350
rect 7803 29339 8111 29348
rect 11230 29404 11538 29413
rect 11230 29402 11236 29404
rect 11292 29402 11316 29404
rect 11372 29402 11396 29404
rect 11452 29402 11476 29404
rect 11532 29402 11538 29404
rect 11292 29350 11294 29402
rect 11474 29350 11476 29402
rect 11230 29348 11236 29350
rect 11292 29348 11316 29350
rect 11372 29348 11396 29350
rect 11452 29348 11476 29350
rect 11532 29348 11538 29350
rect 11230 29339 11538 29348
rect 14657 29404 14965 29413
rect 14657 29402 14663 29404
rect 14719 29402 14743 29404
rect 14799 29402 14823 29404
rect 14879 29402 14903 29404
rect 14959 29402 14965 29404
rect 14719 29350 14721 29402
rect 14901 29350 14903 29402
rect 14657 29348 14663 29350
rect 14719 29348 14743 29350
rect 14799 29348 14823 29350
rect 14879 29348 14903 29350
rect 14959 29348 14965 29350
rect 14657 29339 14965 29348
rect 2663 28860 2971 28869
rect 2663 28858 2669 28860
rect 2725 28858 2749 28860
rect 2805 28858 2829 28860
rect 2885 28858 2909 28860
rect 2965 28858 2971 28860
rect 2725 28806 2727 28858
rect 2907 28806 2909 28858
rect 2663 28804 2669 28806
rect 2725 28804 2749 28806
rect 2805 28804 2829 28806
rect 2885 28804 2909 28806
rect 2965 28804 2971 28806
rect 2663 28795 2971 28804
rect 6090 28860 6398 28869
rect 6090 28858 6096 28860
rect 6152 28858 6176 28860
rect 6232 28858 6256 28860
rect 6312 28858 6336 28860
rect 6392 28858 6398 28860
rect 6152 28806 6154 28858
rect 6334 28806 6336 28858
rect 6090 28804 6096 28806
rect 6152 28804 6176 28806
rect 6232 28804 6256 28806
rect 6312 28804 6336 28806
rect 6392 28804 6398 28806
rect 6090 28795 6398 28804
rect 9517 28860 9825 28869
rect 9517 28858 9523 28860
rect 9579 28858 9603 28860
rect 9659 28858 9683 28860
rect 9739 28858 9763 28860
rect 9819 28858 9825 28860
rect 9579 28806 9581 28858
rect 9761 28806 9763 28858
rect 9517 28804 9523 28806
rect 9579 28804 9603 28806
rect 9659 28804 9683 28806
rect 9739 28804 9763 28806
rect 9819 28804 9825 28806
rect 9517 28795 9825 28804
rect 12944 28860 13252 28869
rect 12944 28858 12950 28860
rect 13006 28858 13030 28860
rect 13086 28858 13110 28860
rect 13166 28858 13190 28860
rect 13246 28858 13252 28860
rect 13006 28806 13008 28858
rect 13188 28806 13190 28858
rect 12944 28804 12950 28806
rect 13006 28804 13030 28806
rect 13086 28804 13110 28806
rect 13166 28804 13190 28806
rect 13246 28804 13252 28806
rect 12944 28795 13252 28804
rect 4376 28316 4684 28325
rect 4376 28314 4382 28316
rect 4438 28314 4462 28316
rect 4518 28314 4542 28316
rect 4598 28314 4622 28316
rect 4678 28314 4684 28316
rect 4438 28262 4440 28314
rect 4620 28262 4622 28314
rect 4376 28260 4382 28262
rect 4438 28260 4462 28262
rect 4518 28260 4542 28262
rect 4598 28260 4622 28262
rect 4678 28260 4684 28262
rect 4376 28251 4684 28260
rect 7803 28316 8111 28325
rect 7803 28314 7809 28316
rect 7865 28314 7889 28316
rect 7945 28314 7969 28316
rect 8025 28314 8049 28316
rect 8105 28314 8111 28316
rect 7865 28262 7867 28314
rect 8047 28262 8049 28314
rect 7803 28260 7809 28262
rect 7865 28260 7889 28262
rect 7945 28260 7969 28262
rect 8025 28260 8049 28262
rect 8105 28260 8111 28262
rect 7803 28251 8111 28260
rect 11230 28316 11538 28325
rect 11230 28314 11236 28316
rect 11292 28314 11316 28316
rect 11372 28314 11396 28316
rect 11452 28314 11476 28316
rect 11532 28314 11538 28316
rect 11292 28262 11294 28314
rect 11474 28262 11476 28314
rect 11230 28260 11236 28262
rect 11292 28260 11316 28262
rect 11372 28260 11396 28262
rect 11452 28260 11476 28262
rect 11532 28260 11538 28262
rect 11230 28251 11538 28260
rect 14657 28316 14965 28325
rect 14657 28314 14663 28316
rect 14719 28314 14743 28316
rect 14799 28314 14823 28316
rect 14879 28314 14903 28316
rect 14959 28314 14965 28316
rect 14719 28262 14721 28314
rect 14901 28262 14903 28314
rect 14657 28260 14663 28262
rect 14719 28260 14743 28262
rect 14799 28260 14823 28262
rect 14879 28260 14903 28262
rect 14959 28260 14965 28262
rect 14657 28251 14965 28260
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14476 27849 14504 27950
rect 14462 27840 14518 27849
rect 2663 27772 2971 27781
rect 2663 27770 2669 27772
rect 2725 27770 2749 27772
rect 2805 27770 2829 27772
rect 2885 27770 2909 27772
rect 2965 27770 2971 27772
rect 2725 27718 2727 27770
rect 2907 27718 2909 27770
rect 2663 27716 2669 27718
rect 2725 27716 2749 27718
rect 2805 27716 2829 27718
rect 2885 27716 2909 27718
rect 2965 27716 2971 27718
rect 2663 27707 2971 27716
rect 6090 27772 6398 27781
rect 6090 27770 6096 27772
rect 6152 27770 6176 27772
rect 6232 27770 6256 27772
rect 6312 27770 6336 27772
rect 6392 27770 6398 27772
rect 6152 27718 6154 27770
rect 6334 27718 6336 27770
rect 6090 27716 6096 27718
rect 6152 27716 6176 27718
rect 6232 27716 6256 27718
rect 6312 27716 6336 27718
rect 6392 27716 6398 27718
rect 6090 27707 6398 27716
rect 9517 27772 9825 27781
rect 9517 27770 9523 27772
rect 9579 27770 9603 27772
rect 9659 27770 9683 27772
rect 9739 27770 9763 27772
rect 9819 27770 9825 27772
rect 9579 27718 9581 27770
rect 9761 27718 9763 27770
rect 9517 27716 9523 27718
rect 9579 27716 9603 27718
rect 9659 27716 9683 27718
rect 9739 27716 9763 27718
rect 9819 27716 9825 27718
rect 9517 27707 9825 27716
rect 12944 27772 13252 27781
rect 14462 27775 14518 27784
rect 12944 27770 12950 27772
rect 13006 27770 13030 27772
rect 13086 27770 13110 27772
rect 13166 27770 13190 27772
rect 13246 27770 13252 27772
rect 13006 27718 13008 27770
rect 13188 27718 13190 27770
rect 12944 27716 12950 27718
rect 13006 27716 13030 27718
rect 13086 27716 13110 27718
rect 13166 27716 13190 27718
rect 13246 27716 13252 27718
rect 12944 27707 13252 27716
rect 4376 27228 4684 27237
rect 4376 27226 4382 27228
rect 4438 27226 4462 27228
rect 4518 27226 4542 27228
rect 4598 27226 4622 27228
rect 4678 27226 4684 27228
rect 4438 27174 4440 27226
rect 4620 27174 4622 27226
rect 4376 27172 4382 27174
rect 4438 27172 4462 27174
rect 4518 27172 4542 27174
rect 4598 27172 4622 27174
rect 4678 27172 4684 27174
rect 4376 27163 4684 27172
rect 7803 27228 8111 27237
rect 7803 27226 7809 27228
rect 7865 27226 7889 27228
rect 7945 27226 7969 27228
rect 8025 27226 8049 27228
rect 8105 27226 8111 27228
rect 7865 27174 7867 27226
rect 8047 27174 8049 27226
rect 7803 27172 7809 27174
rect 7865 27172 7889 27174
rect 7945 27172 7969 27174
rect 8025 27172 8049 27174
rect 8105 27172 8111 27174
rect 7803 27163 8111 27172
rect 11230 27228 11538 27237
rect 11230 27226 11236 27228
rect 11292 27226 11316 27228
rect 11372 27226 11396 27228
rect 11452 27226 11476 27228
rect 11532 27226 11538 27228
rect 11292 27174 11294 27226
rect 11474 27174 11476 27226
rect 11230 27172 11236 27174
rect 11292 27172 11316 27174
rect 11372 27172 11396 27174
rect 11452 27172 11476 27174
rect 11532 27172 11538 27174
rect 11230 27163 11538 27172
rect 14657 27228 14965 27237
rect 14657 27226 14663 27228
rect 14719 27226 14743 27228
rect 14799 27226 14823 27228
rect 14879 27226 14903 27228
rect 14959 27226 14965 27228
rect 14719 27174 14721 27226
rect 14901 27174 14903 27226
rect 14657 27172 14663 27174
rect 14719 27172 14743 27174
rect 14799 27172 14823 27174
rect 14879 27172 14903 27174
rect 14959 27172 14965 27174
rect 14657 27163 14965 27172
rect 2663 26684 2971 26693
rect 2663 26682 2669 26684
rect 2725 26682 2749 26684
rect 2805 26682 2829 26684
rect 2885 26682 2909 26684
rect 2965 26682 2971 26684
rect 2725 26630 2727 26682
rect 2907 26630 2909 26682
rect 2663 26628 2669 26630
rect 2725 26628 2749 26630
rect 2805 26628 2829 26630
rect 2885 26628 2909 26630
rect 2965 26628 2971 26630
rect 2663 26619 2971 26628
rect 6090 26684 6398 26693
rect 6090 26682 6096 26684
rect 6152 26682 6176 26684
rect 6232 26682 6256 26684
rect 6312 26682 6336 26684
rect 6392 26682 6398 26684
rect 6152 26630 6154 26682
rect 6334 26630 6336 26682
rect 6090 26628 6096 26630
rect 6152 26628 6176 26630
rect 6232 26628 6256 26630
rect 6312 26628 6336 26630
rect 6392 26628 6398 26630
rect 6090 26619 6398 26628
rect 9517 26684 9825 26693
rect 9517 26682 9523 26684
rect 9579 26682 9603 26684
rect 9659 26682 9683 26684
rect 9739 26682 9763 26684
rect 9819 26682 9825 26684
rect 9579 26630 9581 26682
rect 9761 26630 9763 26682
rect 9517 26628 9523 26630
rect 9579 26628 9603 26630
rect 9659 26628 9683 26630
rect 9739 26628 9763 26630
rect 9819 26628 9825 26630
rect 9517 26619 9825 26628
rect 12944 26684 13252 26693
rect 12944 26682 12950 26684
rect 13006 26682 13030 26684
rect 13086 26682 13110 26684
rect 13166 26682 13190 26684
rect 13246 26682 13252 26684
rect 13006 26630 13008 26682
rect 13188 26630 13190 26682
rect 12944 26628 12950 26630
rect 13006 26628 13030 26630
rect 13086 26628 13110 26630
rect 13166 26628 13190 26630
rect 13246 26628 13252 26630
rect 12944 26619 13252 26628
rect 4376 26140 4684 26149
rect 4376 26138 4382 26140
rect 4438 26138 4462 26140
rect 4518 26138 4542 26140
rect 4598 26138 4622 26140
rect 4678 26138 4684 26140
rect 4438 26086 4440 26138
rect 4620 26086 4622 26138
rect 4376 26084 4382 26086
rect 4438 26084 4462 26086
rect 4518 26084 4542 26086
rect 4598 26084 4622 26086
rect 4678 26084 4684 26086
rect 4376 26075 4684 26084
rect 7803 26140 8111 26149
rect 7803 26138 7809 26140
rect 7865 26138 7889 26140
rect 7945 26138 7969 26140
rect 8025 26138 8049 26140
rect 8105 26138 8111 26140
rect 7865 26086 7867 26138
rect 8047 26086 8049 26138
rect 7803 26084 7809 26086
rect 7865 26084 7889 26086
rect 7945 26084 7969 26086
rect 8025 26084 8049 26086
rect 8105 26084 8111 26086
rect 7803 26075 8111 26084
rect 11230 26140 11538 26149
rect 11230 26138 11236 26140
rect 11292 26138 11316 26140
rect 11372 26138 11396 26140
rect 11452 26138 11476 26140
rect 11532 26138 11538 26140
rect 11292 26086 11294 26138
rect 11474 26086 11476 26138
rect 11230 26084 11236 26086
rect 11292 26084 11316 26086
rect 11372 26084 11396 26086
rect 11452 26084 11476 26086
rect 11532 26084 11538 26086
rect 11230 26075 11538 26084
rect 14657 26140 14965 26149
rect 14657 26138 14663 26140
rect 14719 26138 14743 26140
rect 14799 26138 14823 26140
rect 14879 26138 14903 26140
rect 14959 26138 14965 26140
rect 14719 26086 14721 26138
rect 14901 26086 14903 26138
rect 14657 26084 14663 26086
rect 14719 26084 14743 26086
rect 14799 26084 14823 26086
rect 14879 26084 14903 26086
rect 14959 26084 14965 26086
rect 14657 26075 14965 26084
rect 2663 25596 2971 25605
rect 2663 25594 2669 25596
rect 2725 25594 2749 25596
rect 2805 25594 2829 25596
rect 2885 25594 2909 25596
rect 2965 25594 2971 25596
rect 2725 25542 2727 25594
rect 2907 25542 2909 25594
rect 2663 25540 2669 25542
rect 2725 25540 2749 25542
rect 2805 25540 2829 25542
rect 2885 25540 2909 25542
rect 2965 25540 2971 25542
rect 2663 25531 2971 25540
rect 6090 25596 6398 25605
rect 6090 25594 6096 25596
rect 6152 25594 6176 25596
rect 6232 25594 6256 25596
rect 6312 25594 6336 25596
rect 6392 25594 6398 25596
rect 6152 25542 6154 25594
rect 6334 25542 6336 25594
rect 6090 25540 6096 25542
rect 6152 25540 6176 25542
rect 6232 25540 6256 25542
rect 6312 25540 6336 25542
rect 6392 25540 6398 25542
rect 6090 25531 6398 25540
rect 9517 25596 9825 25605
rect 9517 25594 9523 25596
rect 9579 25594 9603 25596
rect 9659 25594 9683 25596
rect 9739 25594 9763 25596
rect 9819 25594 9825 25596
rect 9579 25542 9581 25594
rect 9761 25542 9763 25594
rect 9517 25540 9523 25542
rect 9579 25540 9603 25542
rect 9659 25540 9683 25542
rect 9739 25540 9763 25542
rect 9819 25540 9825 25542
rect 9517 25531 9825 25540
rect 12944 25596 13252 25605
rect 12944 25594 12950 25596
rect 13006 25594 13030 25596
rect 13086 25594 13110 25596
rect 13166 25594 13190 25596
rect 13246 25594 13252 25596
rect 13006 25542 13008 25594
rect 13188 25542 13190 25594
rect 12944 25540 12950 25542
rect 13006 25540 13030 25542
rect 13086 25540 13110 25542
rect 13166 25540 13190 25542
rect 13246 25540 13252 25542
rect 12944 25531 13252 25540
rect 4376 25052 4684 25061
rect 4376 25050 4382 25052
rect 4438 25050 4462 25052
rect 4518 25050 4542 25052
rect 4598 25050 4622 25052
rect 4678 25050 4684 25052
rect 4438 24998 4440 25050
rect 4620 24998 4622 25050
rect 4376 24996 4382 24998
rect 4438 24996 4462 24998
rect 4518 24996 4542 24998
rect 4598 24996 4622 24998
rect 4678 24996 4684 24998
rect 4376 24987 4684 24996
rect 7803 25052 8111 25061
rect 7803 25050 7809 25052
rect 7865 25050 7889 25052
rect 7945 25050 7969 25052
rect 8025 25050 8049 25052
rect 8105 25050 8111 25052
rect 7865 24998 7867 25050
rect 8047 24998 8049 25050
rect 7803 24996 7809 24998
rect 7865 24996 7889 24998
rect 7945 24996 7969 24998
rect 8025 24996 8049 24998
rect 8105 24996 8111 24998
rect 7803 24987 8111 24996
rect 11230 25052 11538 25061
rect 11230 25050 11236 25052
rect 11292 25050 11316 25052
rect 11372 25050 11396 25052
rect 11452 25050 11476 25052
rect 11532 25050 11538 25052
rect 11292 24998 11294 25050
rect 11474 24998 11476 25050
rect 11230 24996 11236 24998
rect 11292 24996 11316 24998
rect 11372 24996 11396 24998
rect 11452 24996 11476 24998
rect 11532 24996 11538 24998
rect 11230 24987 11538 24996
rect 14657 25052 14965 25061
rect 14657 25050 14663 25052
rect 14719 25050 14743 25052
rect 14799 25050 14823 25052
rect 14879 25050 14903 25052
rect 14959 25050 14965 25052
rect 14719 24998 14721 25050
rect 14901 24998 14903 25050
rect 14657 24996 14663 24998
rect 14719 24996 14743 24998
rect 14799 24996 14823 24998
rect 14879 24996 14903 24998
rect 14959 24996 14965 24998
rect 14657 24987 14965 24996
rect 2663 24508 2971 24517
rect 2663 24506 2669 24508
rect 2725 24506 2749 24508
rect 2805 24506 2829 24508
rect 2885 24506 2909 24508
rect 2965 24506 2971 24508
rect 2725 24454 2727 24506
rect 2907 24454 2909 24506
rect 2663 24452 2669 24454
rect 2725 24452 2749 24454
rect 2805 24452 2829 24454
rect 2885 24452 2909 24454
rect 2965 24452 2971 24454
rect 2663 24443 2971 24452
rect 6090 24508 6398 24517
rect 6090 24506 6096 24508
rect 6152 24506 6176 24508
rect 6232 24506 6256 24508
rect 6312 24506 6336 24508
rect 6392 24506 6398 24508
rect 6152 24454 6154 24506
rect 6334 24454 6336 24506
rect 6090 24452 6096 24454
rect 6152 24452 6176 24454
rect 6232 24452 6256 24454
rect 6312 24452 6336 24454
rect 6392 24452 6398 24454
rect 6090 24443 6398 24452
rect 9517 24508 9825 24517
rect 9517 24506 9523 24508
rect 9579 24506 9603 24508
rect 9659 24506 9683 24508
rect 9739 24506 9763 24508
rect 9819 24506 9825 24508
rect 9579 24454 9581 24506
rect 9761 24454 9763 24506
rect 9517 24452 9523 24454
rect 9579 24452 9603 24454
rect 9659 24452 9683 24454
rect 9739 24452 9763 24454
rect 9819 24452 9825 24454
rect 9517 24443 9825 24452
rect 12944 24508 13252 24517
rect 12944 24506 12950 24508
rect 13006 24506 13030 24508
rect 13086 24506 13110 24508
rect 13166 24506 13190 24508
rect 13246 24506 13252 24508
rect 13006 24454 13008 24506
rect 13188 24454 13190 24506
rect 12944 24452 12950 24454
rect 13006 24452 13030 24454
rect 13086 24452 13110 24454
rect 13166 24452 13190 24454
rect 13246 24452 13252 24454
rect 12944 24443 13252 24452
rect 4376 23964 4684 23973
rect 4376 23962 4382 23964
rect 4438 23962 4462 23964
rect 4518 23962 4542 23964
rect 4598 23962 4622 23964
rect 4678 23962 4684 23964
rect 4438 23910 4440 23962
rect 4620 23910 4622 23962
rect 4376 23908 4382 23910
rect 4438 23908 4462 23910
rect 4518 23908 4542 23910
rect 4598 23908 4622 23910
rect 4678 23908 4684 23910
rect 4376 23899 4684 23908
rect 7803 23964 8111 23973
rect 7803 23962 7809 23964
rect 7865 23962 7889 23964
rect 7945 23962 7969 23964
rect 8025 23962 8049 23964
rect 8105 23962 8111 23964
rect 7865 23910 7867 23962
rect 8047 23910 8049 23962
rect 7803 23908 7809 23910
rect 7865 23908 7889 23910
rect 7945 23908 7969 23910
rect 8025 23908 8049 23910
rect 8105 23908 8111 23910
rect 7803 23899 8111 23908
rect 11230 23964 11538 23973
rect 11230 23962 11236 23964
rect 11292 23962 11316 23964
rect 11372 23962 11396 23964
rect 11452 23962 11476 23964
rect 11532 23962 11538 23964
rect 11292 23910 11294 23962
rect 11474 23910 11476 23962
rect 11230 23908 11236 23910
rect 11292 23908 11316 23910
rect 11372 23908 11396 23910
rect 11452 23908 11476 23910
rect 11532 23908 11538 23910
rect 11230 23899 11538 23908
rect 14657 23964 14965 23973
rect 14657 23962 14663 23964
rect 14719 23962 14743 23964
rect 14799 23962 14823 23964
rect 14879 23962 14903 23964
rect 14959 23962 14965 23964
rect 14719 23910 14721 23962
rect 14901 23910 14903 23962
rect 14657 23908 14663 23910
rect 14719 23908 14743 23910
rect 14799 23908 14823 23910
rect 14879 23908 14903 23910
rect 14959 23908 14965 23910
rect 14657 23899 14965 23908
rect 2663 23420 2971 23429
rect 2663 23418 2669 23420
rect 2725 23418 2749 23420
rect 2805 23418 2829 23420
rect 2885 23418 2909 23420
rect 2965 23418 2971 23420
rect 2725 23366 2727 23418
rect 2907 23366 2909 23418
rect 2663 23364 2669 23366
rect 2725 23364 2749 23366
rect 2805 23364 2829 23366
rect 2885 23364 2909 23366
rect 2965 23364 2971 23366
rect 2663 23355 2971 23364
rect 6090 23420 6398 23429
rect 6090 23418 6096 23420
rect 6152 23418 6176 23420
rect 6232 23418 6256 23420
rect 6312 23418 6336 23420
rect 6392 23418 6398 23420
rect 6152 23366 6154 23418
rect 6334 23366 6336 23418
rect 6090 23364 6096 23366
rect 6152 23364 6176 23366
rect 6232 23364 6256 23366
rect 6312 23364 6336 23366
rect 6392 23364 6398 23366
rect 6090 23355 6398 23364
rect 9517 23420 9825 23429
rect 9517 23418 9523 23420
rect 9579 23418 9603 23420
rect 9659 23418 9683 23420
rect 9739 23418 9763 23420
rect 9819 23418 9825 23420
rect 9579 23366 9581 23418
rect 9761 23366 9763 23418
rect 9517 23364 9523 23366
rect 9579 23364 9603 23366
rect 9659 23364 9683 23366
rect 9739 23364 9763 23366
rect 9819 23364 9825 23366
rect 9517 23355 9825 23364
rect 12944 23420 13252 23429
rect 12944 23418 12950 23420
rect 13006 23418 13030 23420
rect 13086 23418 13110 23420
rect 13166 23418 13190 23420
rect 13246 23418 13252 23420
rect 13006 23366 13008 23418
rect 13188 23366 13190 23418
rect 12944 23364 12950 23366
rect 13006 23364 13030 23366
rect 13086 23364 13110 23366
rect 13166 23364 13190 23366
rect 13246 23364 13252 23366
rect 12944 23355 13252 23364
rect 4376 22876 4684 22885
rect 4376 22874 4382 22876
rect 4438 22874 4462 22876
rect 4518 22874 4542 22876
rect 4598 22874 4622 22876
rect 4678 22874 4684 22876
rect 4438 22822 4440 22874
rect 4620 22822 4622 22874
rect 4376 22820 4382 22822
rect 4438 22820 4462 22822
rect 4518 22820 4542 22822
rect 4598 22820 4622 22822
rect 4678 22820 4684 22822
rect 4376 22811 4684 22820
rect 7803 22876 8111 22885
rect 7803 22874 7809 22876
rect 7865 22874 7889 22876
rect 7945 22874 7969 22876
rect 8025 22874 8049 22876
rect 8105 22874 8111 22876
rect 7865 22822 7867 22874
rect 8047 22822 8049 22874
rect 7803 22820 7809 22822
rect 7865 22820 7889 22822
rect 7945 22820 7969 22822
rect 8025 22820 8049 22822
rect 8105 22820 8111 22822
rect 7803 22811 8111 22820
rect 11230 22876 11538 22885
rect 11230 22874 11236 22876
rect 11292 22874 11316 22876
rect 11372 22874 11396 22876
rect 11452 22874 11476 22876
rect 11532 22874 11538 22876
rect 11292 22822 11294 22874
rect 11474 22822 11476 22874
rect 11230 22820 11236 22822
rect 11292 22820 11316 22822
rect 11372 22820 11396 22822
rect 11452 22820 11476 22822
rect 11532 22820 11538 22822
rect 11230 22811 11538 22820
rect 14657 22876 14965 22885
rect 14657 22874 14663 22876
rect 14719 22874 14743 22876
rect 14799 22874 14823 22876
rect 14879 22874 14903 22876
rect 14959 22874 14965 22876
rect 14719 22822 14721 22874
rect 14901 22822 14903 22874
rect 14657 22820 14663 22822
rect 14719 22820 14743 22822
rect 14799 22820 14823 22822
rect 14879 22820 14903 22822
rect 14959 22820 14965 22822
rect 14657 22811 14965 22820
rect 2663 22332 2971 22341
rect 2663 22330 2669 22332
rect 2725 22330 2749 22332
rect 2805 22330 2829 22332
rect 2885 22330 2909 22332
rect 2965 22330 2971 22332
rect 2725 22278 2727 22330
rect 2907 22278 2909 22330
rect 2663 22276 2669 22278
rect 2725 22276 2749 22278
rect 2805 22276 2829 22278
rect 2885 22276 2909 22278
rect 2965 22276 2971 22278
rect 2663 22267 2971 22276
rect 6090 22332 6398 22341
rect 6090 22330 6096 22332
rect 6152 22330 6176 22332
rect 6232 22330 6256 22332
rect 6312 22330 6336 22332
rect 6392 22330 6398 22332
rect 6152 22278 6154 22330
rect 6334 22278 6336 22330
rect 6090 22276 6096 22278
rect 6152 22276 6176 22278
rect 6232 22276 6256 22278
rect 6312 22276 6336 22278
rect 6392 22276 6398 22278
rect 6090 22267 6398 22276
rect 9517 22332 9825 22341
rect 9517 22330 9523 22332
rect 9579 22330 9603 22332
rect 9659 22330 9683 22332
rect 9739 22330 9763 22332
rect 9819 22330 9825 22332
rect 9579 22278 9581 22330
rect 9761 22278 9763 22330
rect 9517 22276 9523 22278
rect 9579 22276 9603 22278
rect 9659 22276 9683 22278
rect 9739 22276 9763 22278
rect 9819 22276 9825 22278
rect 9517 22267 9825 22276
rect 12944 22332 13252 22341
rect 12944 22330 12950 22332
rect 13006 22330 13030 22332
rect 13086 22330 13110 22332
rect 13166 22330 13190 22332
rect 13246 22330 13252 22332
rect 13006 22278 13008 22330
rect 13188 22278 13190 22330
rect 12944 22276 12950 22278
rect 13006 22276 13030 22278
rect 13086 22276 13110 22278
rect 13166 22276 13190 22278
rect 13246 22276 13252 22278
rect 12944 22267 13252 22276
rect 4376 21788 4684 21797
rect 4376 21786 4382 21788
rect 4438 21786 4462 21788
rect 4518 21786 4542 21788
rect 4598 21786 4622 21788
rect 4678 21786 4684 21788
rect 4438 21734 4440 21786
rect 4620 21734 4622 21786
rect 4376 21732 4382 21734
rect 4438 21732 4462 21734
rect 4518 21732 4542 21734
rect 4598 21732 4622 21734
rect 4678 21732 4684 21734
rect 4376 21723 4684 21732
rect 7803 21788 8111 21797
rect 7803 21786 7809 21788
rect 7865 21786 7889 21788
rect 7945 21786 7969 21788
rect 8025 21786 8049 21788
rect 8105 21786 8111 21788
rect 7865 21734 7867 21786
rect 8047 21734 8049 21786
rect 7803 21732 7809 21734
rect 7865 21732 7889 21734
rect 7945 21732 7969 21734
rect 8025 21732 8049 21734
rect 8105 21732 8111 21734
rect 7803 21723 8111 21732
rect 11230 21788 11538 21797
rect 11230 21786 11236 21788
rect 11292 21786 11316 21788
rect 11372 21786 11396 21788
rect 11452 21786 11476 21788
rect 11532 21786 11538 21788
rect 11292 21734 11294 21786
rect 11474 21734 11476 21786
rect 11230 21732 11236 21734
rect 11292 21732 11316 21734
rect 11372 21732 11396 21734
rect 11452 21732 11476 21734
rect 11532 21732 11538 21734
rect 11230 21723 11538 21732
rect 14657 21788 14965 21797
rect 14657 21786 14663 21788
rect 14719 21786 14743 21788
rect 14799 21786 14823 21788
rect 14879 21786 14903 21788
rect 14959 21786 14965 21788
rect 14719 21734 14721 21786
rect 14901 21734 14903 21786
rect 14657 21732 14663 21734
rect 14719 21732 14743 21734
rect 14799 21732 14823 21734
rect 14879 21732 14903 21734
rect 14959 21732 14965 21734
rect 14657 21723 14965 21732
rect 2663 21244 2971 21253
rect 2663 21242 2669 21244
rect 2725 21242 2749 21244
rect 2805 21242 2829 21244
rect 2885 21242 2909 21244
rect 2965 21242 2971 21244
rect 2725 21190 2727 21242
rect 2907 21190 2909 21242
rect 2663 21188 2669 21190
rect 2725 21188 2749 21190
rect 2805 21188 2829 21190
rect 2885 21188 2909 21190
rect 2965 21188 2971 21190
rect 2663 21179 2971 21188
rect 6090 21244 6398 21253
rect 6090 21242 6096 21244
rect 6152 21242 6176 21244
rect 6232 21242 6256 21244
rect 6312 21242 6336 21244
rect 6392 21242 6398 21244
rect 6152 21190 6154 21242
rect 6334 21190 6336 21242
rect 6090 21188 6096 21190
rect 6152 21188 6176 21190
rect 6232 21188 6256 21190
rect 6312 21188 6336 21190
rect 6392 21188 6398 21190
rect 6090 21179 6398 21188
rect 9517 21244 9825 21253
rect 9517 21242 9523 21244
rect 9579 21242 9603 21244
rect 9659 21242 9683 21244
rect 9739 21242 9763 21244
rect 9819 21242 9825 21244
rect 9579 21190 9581 21242
rect 9761 21190 9763 21242
rect 9517 21188 9523 21190
rect 9579 21188 9603 21190
rect 9659 21188 9683 21190
rect 9739 21188 9763 21190
rect 9819 21188 9825 21190
rect 9517 21179 9825 21188
rect 12944 21244 13252 21253
rect 12944 21242 12950 21244
rect 13006 21242 13030 21244
rect 13086 21242 13110 21244
rect 13166 21242 13190 21244
rect 13246 21242 13252 21244
rect 13006 21190 13008 21242
rect 13188 21190 13190 21242
rect 12944 21188 12950 21190
rect 13006 21188 13030 21190
rect 13086 21188 13110 21190
rect 13166 21188 13190 21190
rect 13246 21188 13252 21190
rect 12944 21179 13252 21188
rect 4376 20700 4684 20709
rect 4376 20698 4382 20700
rect 4438 20698 4462 20700
rect 4518 20698 4542 20700
rect 4598 20698 4622 20700
rect 4678 20698 4684 20700
rect 4438 20646 4440 20698
rect 4620 20646 4622 20698
rect 4376 20644 4382 20646
rect 4438 20644 4462 20646
rect 4518 20644 4542 20646
rect 4598 20644 4622 20646
rect 4678 20644 4684 20646
rect 4376 20635 4684 20644
rect 7803 20700 8111 20709
rect 7803 20698 7809 20700
rect 7865 20698 7889 20700
rect 7945 20698 7969 20700
rect 8025 20698 8049 20700
rect 8105 20698 8111 20700
rect 7865 20646 7867 20698
rect 8047 20646 8049 20698
rect 7803 20644 7809 20646
rect 7865 20644 7889 20646
rect 7945 20644 7969 20646
rect 8025 20644 8049 20646
rect 8105 20644 8111 20646
rect 7803 20635 8111 20644
rect 11230 20700 11538 20709
rect 11230 20698 11236 20700
rect 11292 20698 11316 20700
rect 11372 20698 11396 20700
rect 11452 20698 11476 20700
rect 11532 20698 11538 20700
rect 11292 20646 11294 20698
rect 11474 20646 11476 20698
rect 11230 20644 11236 20646
rect 11292 20644 11316 20646
rect 11372 20644 11396 20646
rect 11452 20644 11476 20646
rect 11532 20644 11538 20646
rect 11230 20635 11538 20644
rect 14657 20700 14965 20709
rect 14657 20698 14663 20700
rect 14719 20698 14743 20700
rect 14799 20698 14823 20700
rect 14879 20698 14903 20700
rect 14959 20698 14965 20700
rect 14719 20646 14721 20698
rect 14901 20646 14903 20698
rect 14657 20644 14663 20646
rect 14719 20644 14743 20646
rect 14799 20644 14823 20646
rect 14879 20644 14903 20646
rect 14959 20644 14965 20646
rect 14657 20635 14965 20644
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 2663 20156 2971 20165
rect 2663 20154 2669 20156
rect 2725 20154 2749 20156
rect 2805 20154 2829 20156
rect 2885 20154 2909 20156
rect 2965 20154 2971 20156
rect 2725 20102 2727 20154
rect 2907 20102 2909 20154
rect 2663 20100 2669 20102
rect 2725 20100 2749 20102
rect 2805 20100 2829 20102
rect 2885 20100 2909 20102
rect 2965 20100 2971 20102
rect 2663 20091 2971 20100
rect 6090 20156 6398 20165
rect 6090 20154 6096 20156
rect 6152 20154 6176 20156
rect 6232 20154 6256 20156
rect 6312 20154 6336 20156
rect 6392 20154 6398 20156
rect 6152 20102 6154 20154
rect 6334 20102 6336 20154
rect 6090 20100 6096 20102
rect 6152 20100 6176 20102
rect 6232 20100 6256 20102
rect 6312 20100 6336 20102
rect 6392 20100 6398 20102
rect 6090 20091 6398 20100
rect 9517 20156 9825 20165
rect 9517 20154 9523 20156
rect 9579 20154 9603 20156
rect 9659 20154 9683 20156
rect 9739 20154 9763 20156
rect 9819 20154 9825 20156
rect 9579 20102 9581 20154
rect 9761 20102 9763 20154
rect 9517 20100 9523 20102
rect 9579 20100 9603 20102
rect 9659 20100 9683 20102
rect 9739 20100 9763 20102
rect 9819 20100 9825 20102
rect 9517 20091 9825 20100
rect 12944 20156 13252 20165
rect 12944 20154 12950 20156
rect 13006 20154 13030 20156
rect 13086 20154 13110 20156
rect 13166 20154 13190 20156
rect 13246 20154 13252 20156
rect 13006 20102 13008 20154
rect 13188 20102 13190 20154
rect 12944 20100 12950 20102
rect 13006 20100 13030 20102
rect 13086 20100 13110 20102
rect 13166 20100 13190 20102
rect 13246 20100 13252 20102
rect 12944 20091 13252 20100
rect 14476 19961 14504 20334
rect 14462 19952 14518 19961
rect 14462 19887 14518 19896
rect 4376 19612 4684 19621
rect 4376 19610 4382 19612
rect 4438 19610 4462 19612
rect 4518 19610 4542 19612
rect 4598 19610 4622 19612
rect 4678 19610 4684 19612
rect 4438 19558 4440 19610
rect 4620 19558 4622 19610
rect 4376 19556 4382 19558
rect 4438 19556 4462 19558
rect 4518 19556 4542 19558
rect 4598 19556 4622 19558
rect 4678 19556 4684 19558
rect 4376 19547 4684 19556
rect 7803 19612 8111 19621
rect 7803 19610 7809 19612
rect 7865 19610 7889 19612
rect 7945 19610 7969 19612
rect 8025 19610 8049 19612
rect 8105 19610 8111 19612
rect 7865 19558 7867 19610
rect 8047 19558 8049 19610
rect 7803 19556 7809 19558
rect 7865 19556 7889 19558
rect 7945 19556 7969 19558
rect 8025 19556 8049 19558
rect 8105 19556 8111 19558
rect 7803 19547 8111 19556
rect 11230 19612 11538 19621
rect 11230 19610 11236 19612
rect 11292 19610 11316 19612
rect 11372 19610 11396 19612
rect 11452 19610 11476 19612
rect 11532 19610 11538 19612
rect 11292 19558 11294 19610
rect 11474 19558 11476 19610
rect 11230 19556 11236 19558
rect 11292 19556 11316 19558
rect 11372 19556 11396 19558
rect 11452 19556 11476 19558
rect 11532 19556 11538 19558
rect 11230 19547 11538 19556
rect 14657 19612 14965 19621
rect 14657 19610 14663 19612
rect 14719 19610 14743 19612
rect 14799 19610 14823 19612
rect 14879 19610 14903 19612
rect 14959 19610 14965 19612
rect 14719 19558 14721 19610
rect 14901 19558 14903 19610
rect 14657 19556 14663 19558
rect 14719 19556 14743 19558
rect 14799 19556 14823 19558
rect 14879 19556 14903 19558
rect 14959 19556 14965 19558
rect 14657 19547 14965 19556
rect 2663 19068 2971 19077
rect 2663 19066 2669 19068
rect 2725 19066 2749 19068
rect 2805 19066 2829 19068
rect 2885 19066 2909 19068
rect 2965 19066 2971 19068
rect 2725 19014 2727 19066
rect 2907 19014 2909 19066
rect 2663 19012 2669 19014
rect 2725 19012 2749 19014
rect 2805 19012 2829 19014
rect 2885 19012 2909 19014
rect 2965 19012 2971 19014
rect 2663 19003 2971 19012
rect 6090 19068 6398 19077
rect 6090 19066 6096 19068
rect 6152 19066 6176 19068
rect 6232 19066 6256 19068
rect 6312 19066 6336 19068
rect 6392 19066 6398 19068
rect 6152 19014 6154 19066
rect 6334 19014 6336 19066
rect 6090 19012 6096 19014
rect 6152 19012 6176 19014
rect 6232 19012 6256 19014
rect 6312 19012 6336 19014
rect 6392 19012 6398 19014
rect 6090 19003 6398 19012
rect 9517 19068 9825 19077
rect 9517 19066 9523 19068
rect 9579 19066 9603 19068
rect 9659 19066 9683 19068
rect 9739 19066 9763 19068
rect 9819 19066 9825 19068
rect 9579 19014 9581 19066
rect 9761 19014 9763 19066
rect 9517 19012 9523 19014
rect 9579 19012 9603 19014
rect 9659 19012 9683 19014
rect 9739 19012 9763 19014
rect 9819 19012 9825 19014
rect 9517 19003 9825 19012
rect 12944 19068 13252 19077
rect 12944 19066 12950 19068
rect 13006 19066 13030 19068
rect 13086 19066 13110 19068
rect 13166 19066 13190 19068
rect 13246 19066 13252 19068
rect 13006 19014 13008 19066
rect 13188 19014 13190 19066
rect 12944 19012 12950 19014
rect 13006 19012 13030 19014
rect 13086 19012 13110 19014
rect 13166 19012 13190 19014
rect 13246 19012 13252 19014
rect 12944 19003 13252 19012
rect 4376 18524 4684 18533
rect 4376 18522 4382 18524
rect 4438 18522 4462 18524
rect 4518 18522 4542 18524
rect 4598 18522 4622 18524
rect 4678 18522 4684 18524
rect 4438 18470 4440 18522
rect 4620 18470 4622 18522
rect 4376 18468 4382 18470
rect 4438 18468 4462 18470
rect 4518 18468 4542 18470
rect 4598 18468 4622 18470
rect 4678 18468 4684 18470
rect 4376 18459 4684 18468
rect 7803 18524 8111 18533
rect 7803 18522 7809 18524
rect 7865 18522 7889 18524
rect 7945 18522 7969 18524
rect 8025 18522 8049 18524
rect 8105 18522 8111 18524
rect 7865 18470 7867 18522
rect 8047 18470 8049 18522
rect 7803 18468 7809 18470
rect 7865 18468 7889 18470
rect 7945 18468 7969 18470
rect 8025 18468 8049 18470
rect 8105 18468 8111 18470
rect 7803 18459 8111 18468
rect 11230 18524 11538 18533
rect 11230 18522 11236 18524
rect 11292 18522 11316 18524
rect 11372 18522 11396 18524
rect 11452 18522 11476 18524
rect 11532 18522 11538 18524
rect 11292 18470 11294 18522
rect 11474 18470 11476 18522
rect 11230 18468 11236 18470
rect 11292 18468 11316 18470
rect 11372 18468 11396 18470
rect 11452 18468 11476 18470
rect 11532 18468 11538 18470
rect 11230 18459 11538 18468
rect 14657 18524 14965 18533
rect 14657 18522 14663 18524
rect 14719 18522 14743 18524
rect 14799 18522 14823 18524
rect 14879 18522 14903 18524
rect 14959 18522 14965 18524
rect 14719 18470 14721 18522
rect 14901 18470 14903 18522
rect 14657 18468 14663 18470
rect 14719 18468 14743 18470
rect 14799 18468 14823 18470
rect 14879 18468 14903 18470
rect 14959 18468 14965 18470
rect 14657 18459 14965 18468
rect 2663 17980 2971 17989
rect 2663 17978 2669 17980
rect 2725 17978 2749 17980
rect 2805 17978 2829 17980
rect 2885 17978 2909 17980
rect 2965 17978 2971 17980
rect 2725 17926 2727 17978
rect 2907 17926 2909 17978
rect 2663 17924 2669 17926
rect 2725 17924 2749 17926
rect 2805 17924 2829 17926
rect 2885 17924 2909 17926
rect 2965 17924 2971 17926
rect 2663 17915 2971 17924
rect 6090 17980 6398 17989
rect 6090 17978 6096 17980
rect 6152 17978 6176 17980
rect 6232 17978 6256 17980
rect 6312 17978 6336 17980
rect 6392 17978 6398 17980
rect 6152 17926 6154 17978
rect 6334 17926 6336 17978
rect 6090 17924 6096 17926
rect 6152 17924 6176 17926
rect 6232 17924 6256 17926
rect 6312 17924 6336 17926
rect 6392 17924 6398 17926
rect 6090 17915 6398 17924
rect 9517 17980 9825 17989
rect 9517 17978 9523 17980
rect 9579 17978 9603 17980
rect 9659 17978 9683 17980
rect 9739 17978 9763 17980
rect 9819 17978 9825 17980
rect 9579 17926 9581 17978
rect 9761 17926 9763 17978
rect 9517 17924 9523 17926
rect 9579 17924 9603 17926
rect 9659 17924 9683 17926
rect 9739 17924 9763 17926
rect 9819 17924 9825 17926
rect 9517 17915 9825 17924
rect 12944 17980 13252 17989
rect 12944 17978 12950 17980
rect 13006 17978 13030 17980
rect 13086 17978 13110 17980
rect 13166 17978 13190 17980
rect 13246 17978 13252 17980
rect 13006 17926 13008 17978
rect 13188 17926 13190 17978
rect 12944 17924 12950 17926
rect 13006 17924 13030 17926
rect 13086 17924 13110 17926
rect 13166 17924 13190 17926
rect 13246 17924 13252 17926
rect 12944 17915 13252 17924
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 14462 12200 14518 12209
rect 14462 12135 14464 12144
rect 14516 12135 14518 12144
rect 14464 12106 14516 12112
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 14476 4185 14504 4422
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14462 4176 14518 4185
rect 14462 4111 14518 4120
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
<< via2 >>
rect 4382 45722 4438 45724
rect 4462 45722 4518 45724
rect 4542 45722 4598 45724
rect 4622 45722 4678 45724
rect 4382 45670 4428 45722
rect 4428 45670 4438 45722
rect 4462 45670 4492 45722
rect 4492 45670 4504 45722
rect 4504 45670 4518 45722
rect 4542 45670 4556 45722
rect 4556 45670 4568 45722
rect 4568 45670 4598 45722
rect 4622 45670 4632 45722
rect 4632 45670 4678 45722
rect 4382 45668 4438 45670
rect 4462 45668 4518 45670
rect 4542 45668 4598 45670
rect 4622 45668 4678 45670
rect 7809 45722 7865 45724
rect 7889 45722 7945 45724
rect 7969 45722 8025 45724
rect 8049 45722 8105 45724
rect 7809 45670 7855 45722
rect 7855 45670 7865 45722
rect 7889 45670 7919 45722
rect 7919 45670 7931 45722
rect 7931 45670 7945 45722
rect 7969 45670 7983 45722
rect 7983 45670 7995 45722
rect 7995 45670 8025 45722
rect 8049 45670 8059 45722
rect 8059 45670 8105 45722
rect 7809 45668 7865 45670
rect 7889 45668 7945 45670
rect 7969 45668 8025 45670
rect 8049 45668 8105 45670
rect 11236 45722 11292 45724
rect 11316 45722 11372 45724
rect 11396 45722 11452 45724
rect 11476 45722 11532 45724
rect 11236 45670 11282 45722
rect 11282 45670 11292 45722
rect 11316 45670 11346 45722
rect 11346 45670 11358 45722
rect 11358 45670 11372 45722
rect 11396 45670 11410 45722
rect 11410 45670 11422 45722
rect 11422 45670 11452 45722
rect 11476 45670 11486 45722
rect 11486 45670 11532 45722
rect 11236 45668 11292 45670
rect 11316 45668 11372 45670
rect 11396 45668 11452 45670
rect 11476 45668 11532 45670
rect 14663 45722 14719 45724
rect 14743 45722 14799 45724
rect 14823 45722 14879 45724
rect 14903 45722 14959 45724
rect 14663 45670 14709 45722
rect 14709 45670 14719 45722
rect 14743 45670 14773 45722
rect 14773 45670 14785 45722
rect 14785 45670 14799 45722
rect 14823 45670 14837 45722
rect 14837 45670 14849 45722
rect 14849 45670 14879 45722
rect 14903 45670 14913 45722
rect 14913 45670 14959 45722
rect 14663 45668 14719 45670
rect 14743 45668 14799 45670
rect 14823 45668 14879 45670
rect 14903 45668 14959 45670
rect 2669 45178 2725 45180
rect 2749 45178 2805 45180
rect 2829 45178 2885 45180
rect 2909 45178 2965 45180
rect 2669 45126 2715 45178
rect 2715 45126 2725 45178
rect 2749 45126 2779 45178
rect 2779 45126 2791 45178
rect 2791 45126 2805 45178
rect 2829 45126 2843 45178
rect 2843 45126 2855 45178
rect 2855 45126 2885 45178
rect 2909 45126 2919 45178
rect 2919 45126 2965 45178
rect 2669 45124 2725 45126
rect 2749 45124 2805 45126
rect 2829 45124 2885 45126
rect 2909 45124 2965 45126
rect 6096 45178 6152 45180
rect 6176 45178 6232 45180
rect 6256 45178 6312 45180
rect 6336 45178 6392 45180
rect 6096 45126 6142 45178
rect 6142 45126 6152 45178
rect 6176 45126 6206 45178
rect 6206 45126 6218 45178
rect 6218 45126 6232 45178
rect 6256 45126 6270 45178
rect 6270 45126 6282 45178
rect 6282 45126 6312 45178
rect 6336 45126 6346 45178
rect 6346 45126 6392 45178
rect 6096 45124 6152 45126
rect 6176 45124 6232 45126
rect 6256 45124 6312 45126
rect 6336 45124 6392 45126
rect 9523 45178 9579 45180
rect 9603 45178 9659 45180
rect 9683 45178 9739 45180
rect 9763 45178 9819 45180
rect 9523 45126 9569 45178
rect 9569 45126 9579 45178
rect 9603 45126 9633 45178
rect 9633 45126 9645 45178
rect 9645 45126 9659 45178
rect 9683 45126 9697 45178
rect 9697 45126 9709 45178
rect 9709 45126 9739 45178
rect 9763 45126 9773 45178
rect 9773 45126 9819 45178
rect 9523 45124 9579 45126
rect 9603 45124 9659 45126
rect 9683 45124 9739 45126
rect 9763 45124 9819 45126
rect 12950 45178 13006 45180
rect 13030 45178 13086 45180
rect 13110 45178 13166 45180
rect 13190 45178 13246 45180
rect 12950 45126 12996 45178
rect 12996 45126 13006 45178
rect 13030 45126 13060 45178
rect 13060 45126 13072 45178
rect 13072 45126 13086 45178
rect 13110 45126 13124 45178
rect 13124 45126 13136 45178
rect 13136 45126 13166 45178
rect 13190 45126 13200 45178
rect 13200 45126 13246 45178
rect 12950 45124 13006 45126
rect 13030 45124 13086 45126
rect 13110 45124 13166 45126
rect 13190 45124 13246 45126
rect 4382 44634 4438 44636
rect 4462 44634 4518 44636
rect 4542 44634 4598 44636
rect 4622 44634 4678 44636
rect 4382 44582 4428 44634
rect 4428 44582 4438 44634
rect 4462 44582 4492 44634
rect 4492 44582 4504 44634
rect 4504 44582 4518 44634
rect 4542 44582 4556 44634
rect 4556 44582 4568 44634
rect 4568 44582 4598 44634
rect 4622 44582 4632 44634
rect 4632 44582 4678 44634
rect 4382 44580 4438 44582
rect 4462 44580 4518 44582
rect 4542 44580 4598 44582
rect 4622 44580 4678 44582
rect 7809 44634 7865 44636
rect 7889 44634 7945 44636
rect 7969 44634 8025 44636
rect 8049 44634 8105 44636
rect 7809 44582 7855 44634
rect 7855 44582 7865 44634
rect 7889 44582 7919 44634
rect 7919 44582 7931 44634
rect 7931 44582 7945 44634
rect 7969 44582 7983 44634
rect 7983 44582 7995 44634
rect 7995 44582 8025 44634
rect 8049 44582 8059 44634
rect 8059 44582 8105 44634
rect 7809 44580 7865 44582
rect 7889 44580 7945 44582
rect 7969 44580 8025 44582
rect 8049 44580 8105 44582
rect 11236 44634 11292 44636
rect 11316 44634 11372 44636
rect 11396 44634 11452 44636
rect 11476 44634 11532 44636
rect 11236 44582 11282 44634
rect 11282 44582 11292 44634
rect 11316 44582 11346 44634
rect 11346 44582 11358 44634
rect 11358 44582 11372 44634
rect 11396 44582 11410 44634
rect 11410 44582 11422 44634
rect 11422 44582 11452 44634
rect 11476 44582 11486 44634
rect 11486 44582 11532 44634
rect 11236 44580 11292 44582
rect 11316 44580 11372 44582
rect 11396 44580 11452 44582
rect 11476 44580 11532 44582
rect 14663 44634 14719 44636
rect 14743 44634 14799 44636
rect 14823 44634 14879 44636
rect 14903 44634 14959 44636
rect 14663 44582 14709 44634
rect 14709 44582 14719 44634
rect 14743 44582 14773 44634
rect 14773 44582 14785 44634
rect 14785 44582 14799 44634
rect 14823 44582 14837 44634
rect 14837 44582 14849 44634
rect 14849 44582 14879 44634
rect 14903 44582 14913 44634
rect 14913 44582 14959 44634
rect 14663 44580 14719 44582
rect 14743 44580 14799 44582
rect 14823 44580 14879 44582
rect 14903 44580 14959 44582
rect 2669 44090 2725 44092
rect 2749 44090 2805 44092
rect 2829 44090 2885 44092
rect 2909 44090 2965 44092
rect 2669 44038 2715 44090
rect 2715 44038 2725 44090
rect 2749 44038 2779 44090
rect 2779 44038 2791 44090
rect 2791 44038 2805 44090
rect 2829 44038 2843 44090
rect 2843 44038 2855 44090
rect 2855 44038 2885 44090
rect 2909 44038 2919 44090
rect 2919 44038 2965 44090
rect 2669 44036 2725 44038
rect 2749 44036 2805 44038
rect 2829 44036 2885 44038
rect 2909 44036 2965 44038
rect 6096 44090 6152 44092
rect 6176 44090 6232 44092
rect 6256 44090 6312 44092
rect 6336 44090 6392 44092
rect 6096 44038 6142 44090
rect 6142 44038 6152 44090
rect 6176 44038 6206 44090
rect 6206 44038 6218 44090
rect 6218 44038 6232 44090
rect 6256 44038 6270 44090
rect 6270 44038 6282 44090
rect 6282 44038 6312 44090
rect 6336 44038 6346 44090
rect 6346 44038 6392 44090
rect 6096 44036 6152 44038
rect 6176 44036 6232 44038
rect 6256 44036 6312 44038
rect 6336 44036 6392 44038
rect 9523 44090 9579 44092
rect 9603 44090 9659 44092
rect 9683 44090 9739 44092
rect 9763 44090 9819 44092
rect 9523 44038 9569 44090
rect 9569 44038 9579 44090
rect 9603 44038 9633 44090
rect 9633 44038 9645 44090
rect 9645 44038 9659 44090
rect 9683 44038 9697 44090
rect 9697 44038 9709 44090
rect 9709 44038 9739 44090
rect 9763 44038 9773 44090
rect 9773 44038 9819 44090
rect 9523 44036 9579 44038
rect 9603 44036 9659 44038
rect 9683 44036 9739 44038
rect 9763 44036 9819 44038
rect 12950 44090 13006 44092
rect 13030 44090 13086 44092
rect 13110 44090 13166 44092
rect 13190 44090 13246 44092
rect 12950 44038 12996 44090
rect 12996 44038 13006 44090
rect 13030 44038 13060 44090
rect 13060 44038 13072 44090
rect 13072 44038 13086 44090
rect 13110 44038 13124 44090
rect 13124 44038 13136 44090
rect 13136 44038 13166 44090
rect 13190 44038 13200 44090
rect 13200 44038 13246 44090
rect 12950 44036 13006 44038
rect 13030 44036 13086 44038
rect 13110 44036 13166 44038
rect 13190 44036 13246 44038
rect 14462 43716 14518 43752
rect 14462 43696 14464 43716
rect 14464 43696 14516 43716
rect 14516 43696 14518 43716
rect 4382 43546 4438 43548
rect 4462 43546 4518 43548
rect 4542 43546 4598 43548
rect 4622 43546 4678 43548
rect 4382 43494 4428 43546
rect 4428 43494 4438 43546
rect 4462 43494 4492 43546
rect 4492 43494 4504 43546
rect 4504 43494 4518 43546
rect 4542 43494 4556 43546
rect 4556 43494 4568 43546
rect 4568 43494 4598 43546
rect 4622 43494 4632 43546
rect 4632 43494 4678 43546
rect 4382 43492 4438 43494
rect 4462 43492 4518 43494
rect 4542 43492 4598 43494
rect 4622 43492 4678 43494
rect 7809 43546 7865 43548
rect 7889 43546 7945 43548
rect 7969 43546 8025 43548
rect 8049 43546 8105 43548
rect 7809 43494 7855 43546
rect 7855 43494 7865 43546
rect 7889 43494 7919 43546
rect 7919 43494 7931 43546
rect 7931 43494 7945 43546
rect 7969 43494 7983 43546
rect 7983 43494 7995 43546
rect 7995 43494 8025 43546
rect 8049 43494 8059 43546
rect 8059 43494 8105 43546
rect 7809 43492 7865 43494
rect 7889 43492 7945 43494
rect 7969 43492 8025 43494
rect 8049 43492 8105 43494
rect 11236 43546 11292 43548
rect 11316 43546 11372 43548
rect 11396 43546 11452 43548
rect 11476 43546 11532 43548
rect 11236 43494 11282 43546
rect 11282 43494 11292 43546
rect 11316 43494 11346 43546
rect 11346 43494 11358 43546
rect 11358 43494 11372 43546
rect 11396 43494 11410 43546
rect 11410 43494 11422 43546
rect 11422 43494 11452 43546
rect 11476 43494 11486 43546
rect 11486 43494 11532 43546
rect 11236 43492 11292 43494
rect 11316 43492 11372 43494
rect 11396 43492 11452 43494
rect 11476 43492 11532 43494
rect 14663 43546 14719 43548
rect 14743 43546 14799 43548
rect 14823 43546 14879 43548
rect 14903 43546 14959 43548
rect 14663 43494 14709 43546
rect 14709 43494 14719 43546
rect 14743 43494 14773 43546
rect 14773 43494 14785 43546
rect 14785 43494 14799 43546
rect 14823 43494 14837 43546
rect 14837 43494 14849 43546
rect 14849 43494 14879 43546
rect 14903 43494 14913 43546
rect 14913 43494 14959 43546
rect 14663 43492 14719 43494
rect 14743 43492 14799 43494
rect 14823 43492 14879 43494
rect 14903 43492 14959 43494
rect 2669 43002 2725 43004
rect 2749 43002 2805 43004
rect 2829 43002 2885 43004
rect 2909 43002 2965 43004
rect 2669 42950 2715 43002
rect 2715 42950 2725 43002
rect 2749 42950 2779 43002
rect 2779 42950 2791 43002
rect 2791 42950 2805 43002
rect 2829 42950 2843 43002
rect 2843 42950 2855 43002
rect 2855 42950 2885 43002
rect 2909 42950 2919 43002
rect 2919 42950 2965 43002
rect 2669 42948 2725 42950
rect 2749 42948 2805 42950
rect 2829 42948 2885 42950
rect 2909 42948 2965 42950
rect 6096 43002 6152 43004
rect 6176 43002 6232 43004
rect 6256 43002 6312 43004
rect 6336 43002 6392 43004
rect 6096 42950 6142 43002
rect 6142 42950 6152 43002
rect 6176 42950 6206 43002
rect 6206 42950 6218 43002
rect 6218 42950 6232 43002
rect 6256 42950 6270 43002
rect 6270 42950 6282 43002
rect 6282 42950 6312 43002
rect 6336 42950 6346 43002
rect 6346 42950 6392 43002
rect 6096 42948 6152 42950
rect 6176 42948 6232 42950
rect 6256 42948 6312 42950
rect 6336 42948 6392 42950
rect 9523 43002 9579 43004
rect 9603 43002 9659 43004
rect 9683 43002 9739 43004
rect 9763 43002 9819 43004
rect 9523 42950 9569 43002
rect 9569 42950 9579 43002
rect 9603 42950 9633 43002
rect 9633 42950 9645 43002
rect 9645 42950 9659 43002
rect 9683 42950 9697 43002
rect 9697 42950 9709 43002
rect 9709 42950 9739 43002
rect 9763 42950 9773 43002
rect 9773 42950 9819 43002
rect 9523 42948 9579 42950
rect 9603 42948 9659 42950
rect 9683 42948 9739 42950
rect 9763 42948 9819 42950
rect 12950 43002 13006 43004
rect 13030 43002 13086 43004
rect 13110 43002 13166 43004
rect 13190 43002 13246 43004
rect 12950 42950 12996 43002
rect 12996 42950 13006 43002
rect 13030 42950 13060 43002
rect 13060 42950 13072 43002
rect 13072 42950 13086 43002
rect 13110 42950 13124 43002
rect 13124 42950 13136 43002
rect 13136 42950 13166 43002
rect 13190 42950 13200 43002
rect 13200 42950 13246 43002
rect 12950 42948 13006 42950
rect 13030 42948 13086 42950
rect 13110 42948 13166 42950
rect 13190 42948 13246 42950
rect 4382 42458 4438 42460
rect 4462 42458 4518 42460
rect 4542 42458 4598 42460
rect 4622 42458 4678 42460
rect 4382 42406 4428 42458
rect 4428 42406 4438 42458
rect 4462 42406 4492 42458
rect 4492 42406 4504 42458
rect 4504 42406 4518 42458
rect 4542 42406 4556 42458
rect 4556 42406 4568 42458
rect 4568 42406 4598 42458
rect 4622 42406 4632 42458
rect 4632 42406 4678 42458
rect 4382 42404 4438 42406
rect 4462 42404 4518 42406
rect 4542 42404 4598 42406
rect 4622 42404 4678 42406
rect 7809 42458 7865 42460
rect 7889 42458 7945 42460
rect 7969 42458 8025 42460
rect 8049 42458 8105 42460
rect 7809 42406 7855 42458
rect 7855 42406 7865 42458
rect 7889 42406 7919 42458
rect 7919 42406 7931 42458
rect 7931 42406 7945 42458
rect 7969 42406 7983 42458
rect 7983 42406 7995 42458
rect 7995 42406 8025 42458
rect 8049 42406 8059 42458
rect 8059 42406 8105 42458
rect 7809 42404 7865 42406
rect 7889 42404 7945 42406
rect 7969 42404 8025 42406
rect 8049 42404 8105 42406
rect 11236 42458 11292 42460
rect 11316 42458 11372 42460
rect 11396 42458 11452 42460
rect 11476 42458 11532 42460
rect 11236 42406 11282 42458
rect 11282 42406 11292 42458
rect 11316 42406 11346 42458
rect 11346 42406 11358 42458
rect 11358 42406 11372 42458
rect 11396 42406 11410 42458
rect 11410 42406 11422 42458
rect 11422 42406 11452 42458
rect 11476 42406 11486 42458
rect 11486 42406 11532 42458
rect 11236 42404 11292 42406
rect 11316 42404 11372 42406
rect 11396 42404 11452 42406
rect 11476 42404 11532 42406
rect 14663 42458 14719 42460
rect 14743 42458 14799 42460
rect 14823 42458 14879 42460
rect 14903 42458 14959 42460
rect 14663 42406 14709 42458
rect 14709 42406 14719 42458
rect 14743 42406 14773 42458
rect 14773 42406 14785 42458
rect 14785 42406 14799 42458
rect 14823 42406 14837 42458
rect 14837 42406 14849 42458
rect 14849 42406 14879 42458
rect 14903 42406 14913 42458
rect 14913 42406 14959 42458
rect 14663 42404 14719 42406
rect 14743 42404 14799 42406
rect 14823 42404 14879 42406
rect 14903 42404 14959 42406
rect 2669 41914 2725 41916
rect 2749 41914 2805 41916
rect 2829 41914 2885 41916
rect 2909 41914 2965 41916
rect 2669 41862 2715 41914
rect 2715 41862 2725 41914
rect 2749 41862 2779 41914
rect 2779 41862 2791 41914
rect 2791 41862 2805 41914
rect 2829 41862 2843 41914
rect 2843 41862 2855 41914
rect 2855 41862 2885 41914
rect 2909 41862 2919 41914
rect 2919 41862 2965 41914
rect 2669 41860 2725 41862
rect 2749 41860 2805 41862
rect 2829 41860 2885 41862
rect 2909 41860 2965 41862
rect 6096 41914 6152 41916
rect 6176 41914 6232 41916
rect 6256 41914 6312 41916
rect 6336 41914 6392 41916
rect 6096 41862 6142 41914
rect 6142 41862 6152 41914
rect 6176 41862 6206 41914
rect 6206 41862 6218 41914
rect 6218 41862 6232 41914
rect 6256 41862 6270 41914
rect 6270 41862 6282 41914
rect 6282 41862 6312 41914
rect 6336 41862 6346 41914
rect 6346 41862 6392 41914
rect 6096 41860 6152 41862
rect 6176 41860 6232 41862
rect 6256 41860 6312 41862
rect 6336 41860 6392 41862
rect 9523 41914 9579 41916
rect 9603 41914 9659 41916
rect 9683 41914 9739 41916
rect 9763 41914 9819 41916
rect 9523 41862 9569 41914
rect 9569 41862 9579 41914
rect 9603 41862 9633 41914
rect 9633 41862 9645 41914
rect 9645 41862 9659 41914
rect 9683 41862 9697 41914
rect 9697 41862 9709 41914
rect 9709 41862 9739 41914
rect 9763 41862 9773 41914
rect 9773 41862 9819 41914
rect 9523 41860 9579 41862
rect 9603 41860 9659 41862
rect 9683 41860 9739 41862
rect 9763 41860 9819 41862
rect 12950 41914 13006 41916
rect 13030 41914 13086 41916
rect 13110 41914 13166 41916
rect 13190 41914 13246 41916
rect 12950 41862 12996 41914
rect 12996 41862 13006 41914
rect 13030 41862 13060 41914
rect 13060 41862 13072 41914
rect 13072 41862 13086 41914
rect 13110 41862 13124 41914
rect 13124 41862 13136 41914
rect 13136 41862 13166 41914
rect 13190 41862 13200 41914
rect 13200 41862 13246 41914
rect 12950 41860 13006 41862
rect 13030 41860 13086 41862
rect 13110 41860 13166 41862
rect 13190 41860 13246 41862
rect 4382 41370 4438 41372
rect 4462 41370 4518 41372
rect 4542 41370 4598 41372
rect 4622 41370 4678 41372
rect 4382 41318 4428 41370
rect 4428 41318 4438 41370
rect 4462 41318 4492 41370
rect 4492 41318 4504 41370
rect 4504 41318 4518 41370
rect 4542 41318 4556 41370
rect 4556 41318 4568 41370
rect 4568 41318 4598 41370
rect 4622 41318 4632 41370
rect 4632 41318 4678 41370
rect 4382 41316 4438 41318
rect 4462 41316 4518 41318
rect 4542 41316 4598 41318
rect 4622 41316 4678 41318
rect 7809 41370 7865 41372
rect 7889 41370 7945 41372
rect 7969 41370 8025 41372
rect 8049 41370 8105 41372
rect 7809 41318 7855 41370
rect 7855 41318 7865 41370
rect 7889 41318 7919 41370
rect 7919 41318 7931 41370
rect 7931 41318 7945 41370
rect 7969 41318 7983 41370
rect 7983 41318 7995 41370
rect 7995 41318 8025 41370
rect 8049 41318 8059 41370
rect 8059 41318 8105 41370
rect 7809 41316 7865 41318
rect 7889 41316 7945 41318
rect 7969 41316 8025 41318
rect 8049 41316 8105 41318
rect 11236 41370 11292 41372
rect 11316 41370 11372 41372
rect 11396 41370 11452 41372
rect 11476 41370 11532 41372
rect 11236 41318 11282 41370
rect 11282 41318 11292 41370
rect 11316 41318 11346 41370
rect 11346 41318 11358 41370
rect 11358 41318 11372 41370
rect 11396 41318 11410 41370
rect 11410 41318 11422 41370
rect 11422 41318 11452 41370
rect 11476 41318 11486 41370
rect 11486 41318 11532 41370
rect 11236 41316 11292 41318
rect 11316 41316 11372 41318
rect 11396 41316 11452 41318
rect 11476 41316 11532 41318
rect 14663 41370 14719 41372
rect 14743 41370 14799 41372
rect 14823 41370 14879 41372
rect 14903 41370 14959 41372
rect 14663 41318 14709 41370
rect 14709 41318 14719 41370
rect 14743 41318 14773 41370
rect 14773 41318 14785 41370
rect 14785 41318 14799 41370
rect 14823 41318 14837 41370
rect 14837 41318 14849 41370
rect 14849 41318 14879 41370
rect 14903 41318 14913 41370
rect 14913 41318 14959 41370
rect 14663 41316 14719 41318
rect 14743 41316 14799 41318
rect 14823 41316 14879 41318
rect 14903 41316 14959 41318
rect 2669 40826 2725 40828
rect 2749 40826 2805 40828
rect 2829 40826 2885 40828
rect 2909 40826 2965 40828
rect 2669 40774 2715 40826
rect 2715 40774 2725 40826
rect 2749 40774 2779 40826
rect 2779 40774 2791 40826
rect 2791 40774 2805 40826
rect 2829 40774 2843 40826
rect 2843 40774 2855 40826
rect 2855 40774 2885 40826
rect 2909 40774 2919 40826
rect 2919 40774 2965 40826
rect 2669 40772 2725 40774
rect 2749 40772 2805 40774
rect 2829 40772 2885 40774
rect 2909 40772 2965 40774
rect 6096 40826 6152 40828
rect 6176 40826 6232 40828
rect 6256 40826 6312 40828
rect 6336 40826 6392 40828
rect 6096 40774 6142 40826
rect 6142 40774 6152 40826
rect 6176 40774 6206 40826
rect 6206 40774 6218 40826
rect 6218 40774 6232 40826
rect 6256 40774 6270 40826
rect 6270 40774 6282 40826
rect 6282 40774 6312 40826
rect 6336 40774 6346 40826
rect 6346 40774 6392 40826
rect 6096 40772 6152 40774
rect 6176 40772 6232 40774
rect 6256 40772 6312 40774
rect 6336 40772 6392 40774
rect 9523 40826 9579 40828
rect 9603 40826 9659 40828
rect 9683 40826 9739 40828
rect 9763 40826 9819 40828
rect 9523 40774 9569 40826
rect 9569 40774 9579 40826
rect 9603 40774 9633 40826
rect 9633 40774 9645 40826
rect 9645 40774 9659 40826
rect 9683 40774 9697 40826
rect 9697 40774 9709 40826
rect 9709 40774 9739 40826
rect 9763 40774 9773 40826
rect 9773 40774 9819 40826
rect 9523 40772 9579 40774
rect 9603 40772 9659 40774
rect 9683 40772 9739 40774
rect 9763 40772 9819 40774
rect 12950 40826 13006 40828
rect 13030 40826 13086 40828
rect 13110 40826 13166 40828
rect 13190 40826 13246 40828
rect 12950 40774 12996 40826
rect 12996 40774 13006 40826
rect 13030 40774 13060 40826
rect 13060 40774 13072 40826
rect 13072 40774 13086 40826
rect 13110 40774 13124 40826
rect 13124 40774 13136 40826
rect 13136 40774 13166 40826
rect 13190 40774 13200 40826
rect 13200 40774 13246 40826
rect 12950 40772 13006 40774
rect 13030 40772 13086 40774
rect 13110 40772 13166 40774
rect 13190 40772 13246 40774
rect 4382 40282 4438 40284
rect 4462 40282 4518 40284
rect 4542 40282 4598 40284
rect 4622 40282 4678 40284
rect 4382 40230 4428 40282
rect 4428 40230 4438 40282
rect 4462 40230 4492 40282
rect 4492 40230 4504 40282
rect 4504 40230 4518 40282
rect 4542 40230 4556 40282
rect 4556 40230 4568 40282
rect 4568 40230 4598 40282
rect 4622 40230 4632 40282
rect 4632 40230 4678 40282
rect 4382 40228 4438 40230
rect 4462 40228 4518 40230
rect 4542 40228 4598 40230
rect 4622 40228 4678 40230
rect 7809 40282 7865 40284
rect 7889 40282 7945 40284
rect 7969 40282 8025 40284
rect 8049 40282 8105 40284
rect 7809 40230 7855 40282
rect 7855 40230 7865 40282
rect 7889 40230 7919 40282
rect 7919 40230 7931 40282
rect 7931 40230 7945 40282
rect 7969 40230 7983 40282
rect 7983 40230 7995 40282
rect 7995 40230 8025 40282
rect 8049 40230 8059 40282
rect 8059 40230 8105 40282
rect 7809 40228 7865 40230
rect 7889 40228 7945 40230
rect 7969 40228 8025 40230
rect 8049 40228 8105 40230
rect 11236 40282 11292 40284
rect 11316 40282 11372 40284
rect 11396 40282 11452 40284
rect 11476 40282 11532 40284
rect 11236 40230 11282 40282
rect 11282 40230 11292 40282
rect 11316 40230 11346 40282
rect 11346 40230 11358 40282
rect 11358 40230 11372 40282
rect 11396 40230 11410 40282
rect 11410 40230 11422 40282
rect 11422 40230 11452 40282
rect 11476 40230 11486 40282
rect 11486 40230 11532 40282
rect 11236 40228 11292 40230
rect 11316 40228 11372 40230
rect 11396 40228 11452 40230
rect 11476 40228 11532 40230
rect 14663 40282 14719 40284
rect 14743 40282 14799 40284
rect 14823 40282 14879 40284
rect 14903 40282 14959 40284
rect 14663 40230 14709 40282
rect 14709 40230 14719 40282
rect 14743 40230 14773 40282
rect 14773 40230 14785 40282
rect 14785 40230 14799 40282
rect 14823 40230 14837 40282
rect 14837 40230 14849 40282
rect 14849 40230 14879 40282
rect 14903 40230 14913 40282
rect 14913 40230 14959 40282
rect 14663 40228 14719 40230
rect 14743 40228 14799 40230
rect 14823 40228 14879 40230
rect 14903 40228 14959 40230
rect 2669 39738 2725 39740
rect 2749 39738 2805 39740
rect 2829 39738 2885 39740
rect 2909 39738 2965 39740
rect 2669 39686 2715 39738
rect 2715 39686 2725 39738
rect 2749 39686 2779 39738
rect 2779 39686 2791 39738
rect 2791 39686 2805 39738
rect 2829 39686 2843 39738
rect 2843 39686 2855 39738
rect 2855 39686 2885 39738
rect 2909 39686 2919 39738
rect 2919 39686 2965 39738
rect 2669 39684 2725 39686
rect 2749 39684 2805 39686
rect 2829 39684 2885 39686
rect 2909 39684 2965 39686
rect 6096 39738 6152 39740
rect 6176 39738 6232 39740
rect 6256 39738 6312 39740
rect 6336 39738 6392 39740
rect 6096 39686 6142 39738
rect 6142 39686 6152 39738
rect 6176 39686 6206 39738
rect 6206 39686 6218 39738
rect 6218 39686 6232 39738
rect 6256 39686 6270 39738
rect 6270 39686 6282 39738
rect 6282 39686 6312 39738
rect 6336 39686 6346 39738
rect 6346 39686 6392 39738
rect 6096 39684 6152 39686
rect 6176 39684 6232 39686
rect 6256 39684 6312 39686
rect 6336 39684 6392 39686
rect 9523 39738 9579 39740
rect 9603 39738 9659 39740
rect 9683 39738 9739 39740
rect 9763 39738 9819 39740
rect 9523 39686 9569 39738
rect 9569 39686 9579 39738
rect 9603 39686 9633 39738
rect 9633 39686 9645 39738
rect 9645 39686 9659 39738
rect 9683 39686 9697 39738
rect 9697 39686 9709 39738
rect 9709 39686 9739 39738
rect 9763 39686 9773 39738
rect 9773 39686 9819 39738
rect 9523 39684 9579 39686
rect 9603 39684 9659 39686
rect 9683 39684 9739 39686
rect 9763 39684 9819 39686
rect 12950 39738 13006 39740
rect 13030 39738 13086 39740
rect 13110 39738 13166 39740
rect 13190 39738 13246 39740
rect 12950 39686 12996 39738
rect 12996 39686 13006 39738
rect 13030 39686 13060 39738
rect 13060 39686 13072 39738
rect 13072 39686 13086 39738
rect 13110 39686 13124 39738
rect 13124 39686 13136 39738
rect 13136 39686 13166 39738
rect 13190 39686 13200 39738
rect 13200 39686 13246 39738
rect 12950 39684 13006 39686
rect 13030 39684 13086 39686
rect 13110 39684 13166 39686
rect 13190 39684 13246 39686
rect 4382 39194 4438 39196
rect 4462 39194 4518 39196
rect 4542 39194 4598 39196
rect 4622 39194 4678 39196
rect 4382 39142 4428 39194
rect 4428 39142 4438 39194
rect 4462 39142 4492 39194
rect 4492 39142 4504 39194
rect 4504 39142 4518 39194
rect 4542 39142 4556 39194
rect 4556 39142 4568 39194
rect 4568 39142 4598 39194
rect 4622 39142 4632 39194
rect 4632 39142 4678 39194
rect 4382 39140 4438 39142
rect 4462 39140 4518 39142
rect 4542 39140 4598 39142
rect 4622 39140 4678 39142
rect 7809 39194 7865 39196
rect 7889 39194 7945 39196
rect 7969 39194 8025 39196
rect 8049 39194 8105 39196
rect 7809 39142 7855 39194
rect 7855 39142 7865 39194
rect 7889 39142 7919 39194
rect 7919 39142 7931 39194
rect 7931 39142 7945 39194
rect 7969 39142 7983 39194
rect 7983 39142 7995 39194
rect 7995 39142 8025 39194
rect 8049 39142 8059 39194
rect 8059 39142 8105 39194
rect 7809 39140 7865 39142
rect 7889 39140 7945 39142
rect 7969 39140 8025 39142
rect 8049 39140 8105 39142
rect 11236 39194 11292 39196
rect 11316 39194 11372 39196
rect 11396 39194 11452 39196
rect 11476 39194 11532 39196
rect 11236 39142 11282 39194
rect 11282 39142 11292 39194
rect 11316 39142 11346 39194
rect 11346 39142 11358 39194
rect 11358 39142 11372 39194
rect 11396 39142 11410 39194
rect 11410 39142 11422 39194
rect 11422 39142 11452 39194
rect 11476 39142 11486 39194
rect 11486 39142 11532 39194
rect 11236 39140 11292 39142
rect 11316 39140 11372 39142
rect 11396 39140 11452 39142
rect 11476 39140 11532 39142
rect 14663 39194 14719 39196
rect 14743 39194 14799 39196
rect 14823 39194 14879 39196
rect 14903 39194 14959 39196
rect 14663 39142 14709 39194
rect 14709 39142 14719 39194
rect 14743 39142 14773 39194
rect 14773 39142 14785 39194
rect 14785 39142 14799 39194
rect 14823 39142 14837 39194
rect 14837 39142 14849 39194
rect 14849 39142 14879 39194
rect 14903 39142 14913 39194
rect 14913 39142 14959 39194
rect 14663 39140 14719 39142
rect 14743 39140 14799 39142
rect 14823 39140 14879 39142
rect 14903 39140 14959 39142
rect 2669 38650 2725 38652
rect 2749 38650 2805 38652
rect 2829 38650 2885 38652
rect 2909 38650 2965 38652
rect 2669 38598 2715 38650
rect 2715 38598 2725 38650
rect 2749 38598 2779 38650
rect 2779 38598 2791 38650
rect 2791 38598 2805 38650
rect 2829 38598 2843 38650
rect 2843 38598 2855 38650
rect 2855 38598 2885 38650
rect 2909 38598 2919 38650
rect 2919 38598 2965 38650
rect 2669 38596 2725 38598
rect 2749 38596 2805 38598
rect 2829 38596 2885 38598
rect 2909 38596 2965 38598
rect 6096 38650 6152 38652
rect 6176 38650 6232 38652
rect 6256 38650 6312 38652
rect 6336 38650 6392 38652
rect 6096 38598 6142 38650
rect 6142 38598 6152 38650
rect 6176 38598 6206 38650
rect 6206 38598 6218 38650
rect 6218 38598 6232 38650
rect 6256 38598 6270 38650
rect 6270 38598 6282 38650
rect 6282 38598 6312 38650
rect 6336 38598 6346 38650
rect 6346 38598 6392 38650
rect 6096 38596 6152 38598
rect 6176 38596 6232 38598
rect 6256 38596 6312 38598
rect 6336 38596 6392 38598
rect 9523 38650 9579 38652
rect 9603 38650 9659 38652
rect 9683 38650 9739 38652
rect 9763 38650 9819 38652
rect 9523 38598 9569 38650
rect 9569 38598 9579 38650
rect 9603 38598 9633 38650
rect 9633 38598 9645 38650
rect 9645 38598 9659 38650
rect 9683 38598 9697 38650
rect 9697 38598 9709 38650
rect 9709 38598 9739 38650
rect 9763 38598 9773 38650
rect 9773 38598 9819 38650
rect 9523 38596 9579 38598
rect 9603 38596 9659 38598
rect 9683 38596 9739 38598
rect 9763 38596 9819 38598
rect 12950 38650 13006 38652
rect 13030 38650 13086 38652
rect 13110 38650 13166 38652
rect 13190 38650 13246 38652
rect 12950 38598 12996 38650
rect 12996 38598 13006 38650
rect 13030 38598 13060 38650
rect 13060 38598 13072 38650
rect 13072 38598 13086 38650
rect 13110 38598 13124 38650
rect 13124 38598 13136 38650
rect 13136 38598 13166 38650
rect 13190 38598 13200 38650
rect 13200 38598 13246 38650
rect 12950 38596 13006 38598
rect 13030 38596 13086 38598
rect 13110 38596 13166 38598
rect 13190 38596 13246 38598
rect 4382 38106 4438 38108
rect 4462 38106 4518 38108
rect 4542 38106 4598 38108
rect 4622 38106 4678 38108
rect 4382 38054 4428 38106
rect 4428 38054 4438 38106
rect 4462 38054 4492 38106
rect 4492 38054 4504 38106
rect 4504 38054 4518 38106
rect 4542 38054 4556 38106
rect 4556 38054 4568 38106
rect 4568 38054 4598 38106
rect 4622 38054 4632 38106
rect 4632 38054 4678 38106
rect 4382 38052 4438 38054
rect 4462 38052 4518 38054
rect 4542 38052 4598 38054
rect 4622 38052 4678 38054
rect 7809 38106 7865 38108
rect 7889 38106 7945 38108
rect 7969 38106 8025 38108
rect 8049 38106 8105 38108
rect 7809 38054 7855 38106
rect 7855 38054 7865 38106
rect 7889 38054 7919 38106
rect 7919 38054 7931 38106
rect 7931 38054 7945 38106
rect 7969 38054 7983 38106
rect 7983 38054 7995 38106
rect 7995 38054 8025 38106
rect 8049 38054 8059 38106
rect 8059 38054 8105 38106
rect 7809 38052 7865 38054
rect 7889 38052 7945 38054
rect 7969 38052 8025 38054
rect 8049 38052 8105 38054
rect 11236 38106 11292 38108
rect 11316 38106 11372 38108
rect 11396 38106 11452 38108
rect 11476 38106 11532 38108
rect 11236 38054 11282 38106
rect 11282 38054 11292 38106
rect 11316 38054 11346 38106
rect 11346 38054 11358 38106
rect 11358 38054 11372 38106
rect 11396 38054 11410 38106
rect 11410 38054 11422 38106
rect 11422 38054 11452 38106
rect 11476 38054 11486 38106
rect 11486 38054 11532 38106
rect 11236 38052 11292 38054
rect 11316 38052 11372 38054
rect 11396 38052 11452 38054
rect 11476 38052 11532 38054
rect 14663 38106 14719 38108
rect 14743 38106 14799 38108
rect 14823 38106 14879 38108
rect 14903 38106 14959 38108
rect 14663 38054 14709 38106
rect 14709 38054 14719 38106
rect 14743 38054 14773 38106
rect 14773 38054 14785 38106
rect 14785 38054 14799 38106
rect 14823 38054 14837 38106
rect 14837 38054 14849 38106
rect 14849 38054 14879 38106
rect 14903 38054 14913 38106
rect 14913 38054 14959 38106
rect 14663 38052 14719 38054
rect 14743 38052 14799 38054
rect 14823 38052 14879 38054
rect 14903 38052 14959 38054
rect 2669 37562 2725 37564
rect 2749 37562 2805 37564
rect 2829 37562 2885 37564
rect 2909 37562 2965 37564
rect 2669 37510 2715 37562
rect 2715 37510 2725 37562
rect 2749 37510 2779 37562
rect 2779 37510 2791 37562
rect 2791 37510 2805 37562
rect 2829 37510 2843 37562
rect 2843 37510 2855 37562
rect 2855 37510 2885 37562
rect 2909 37510 2919 37562
rect 2919 37510 2965 37562
rect 2669 37508 2725 37510
rect 2749 37508 2805 37510
rect 2829 37508 2885 37510
rect 2909 37508 2965 37510
rect 6096 37562 6152 37564
rect 6176 37562 6232 37564
rect 6256 37562 6312 37564
rect 6336 37562 6392 37564
rect 6096 37510 6142 37562
rect 6142 37510 6152 37562
rect 6176 37510 6206 37562
rect 6206 37510 6218 37562
rect 6218 37510 6232 37562
rect 6256 37510 6270 37562
rect 6270 37510 6282 37562
rect 6282 37510 6312 37562
rect 6336 37510 6346 37562
rect 6346 37510 6392 37562
rect 6096 37508 6152 37510
rect 6176 37508 6232 37510
rect 6256 37508 6312 37510
rect 6336 37508 6392 37510
rect 9523 37562 9579 37564
rect 9603 37562 9659 37564
rect 9683 37562 9739 37564
rect 9763 37562 9819 37564
rect 9523 37510 9569 37562
rect 9569 37510 9579 37562
rect 9603 37510 9633 37562
rect 9633 37510 9645 37562
rect 9645 37510 9659 37562
rect 9683 37510 9697 37562
rect 9697 37510 9709 37562
rect 9709 37510 9739 37562
rect 9763 37510 9773 37562
rect 9773 37510 9819 37562
rect 9523 37508 9579 37510
rect 9603 37508 9659 37510
rect 9683 37508 9739 37510
rect 9763 37508 9819 37510
rect 12950 37562 13006 37564
rect 13030 37562 13086 37564
rect 13110 37562 13166 37564
rect 13190 37562 13246 37564
rect 12950 37510 12996 37562
rect 12996 37510 13006 37562
rect 13030 37510 13060 37562
rect 13060 37510 13072 37562
rect 13072 37510 13086 37562
rect 13110 37510 13124 37562
rect 13124 37510 13136 37562
rect 13136 37510 13166 37562
rect 13190 37510 13200 37562
rect 13200 37510 13246 37562
rect 12950 37508 13006 37510
rect 13030 37508 13086 37510
rect 13110 37508 13166 37510
rect 13190 37508 13246 37510
rect 4382 37018 4438 37020
rect 4462 37018 4518 37020
rect 4542 37018 4598 37020
rect 4622 37018 4678 37020
rect 4382 36966 4428 37018
rect 4428 36966 4438 37018
rect 4462 36966 4492 37018
rect 4492 36966 4504 37018
rect 4504 36966 4518 37018
rect 4542 36966 4556 37018
rect 4556 36966 4568 37018
rect 4568 36966 4598 37018
rect 4622 36966 4632 37018
rect 4632 36966 4678 37018
rect 4382 36964 4438 36966
rect 4462 36964 4518 36966
rect 4542 36964 4598 36966
rect 4622 36964 4678 36966
rect 7809 37018 7865 37020
rect 7889 37018 7945 37020
rect 7969 37018 8025 37020
rect 8049 37018 8105 37020
rect 7809 36966 7855 37018
rect 7855 36966 7865 37018
rect 7889 36966 7919 37018
rect 7919 36966 7931 37018
rect 7931 36966 7945 37018
rect 7969 36966 7983 37018
rect 7983 36966 7995 37018
rect 7995 36966 8025 37018
rect 8049 36966 8059 37018
rect 8059 36966 8105 37018
rect 7809 36964 7865 36966
rect 7889 36964 7945 36966
rect 7969 36964 8025 36966
rect 8049 36964 8105 36966
rect 11236 37018 11292 37020
rect 11316 37018 11372 37020
rect 11396 37018 11452 37020
rect 11476 37018 11532 37020
rect 11236 36966 11282 37018
rect 11282 36966 11292 37018
rect 11316 36966 11346 37018
rect 11346 36966 11358 37018
rect 11358 36966 11372 37018
rect 11396 36966 11410 37018
rect 11410 36966 11422 37018
rect 11422 36966 11452 37018
rect 11476 36966 11486 37018
rect 11486 36966 11532 37018
rect 11236 36964 11292 36966
rect 11316 36964 11372 36966
rect 11396 36964 11452 36966
rect 11476 36964 11532 36966
rect 14663 37018 14719 37020
rect 14743 37018 14799 37020
rect 14823 37018 14879 37020
rect 14903 37018 14959 37020
rect 14663 36966 14709 37018
rect 14709 36966 14719 37018
rect 14743 36966 14773 37018
rect 14773 36966 14785 37018
rect 14785 36966 14799 37018
rect 14823 36966 14837 37018
rect 14837 36966 14849 37018
rect 14849 36966 14879 37018
rect 14903 36966 14913 37018
rect 14913 36966 14959 37018
rect 14663 36964 14719 36966
rect 14743 36964 14799 36966
rect 14823 36964 14879 36966
rect 14903 36964 14959 36966
rect 2669 36474 2725 36476
rect 2749 36474 2805 36476
rect 2829 36474 2885 36476
rect 2909 36474 2965 36476
rect 2669 36422 2715 36474
rect 2715 36422 2725 36474
rect 2749 36422 2779 36474
rect 2779 36422 2791 36474
rect 2791 36422 2805 36474
rect 2829 36422 2843 36474
rect 2843 36422 2855 36474
rect 2855 36422 2885 36474
rect 2909 36422 2919 36474
rect 2919 36422 2965 36474
rect 2669 36420 2725 36422
rect 2749 36420 2805 36422
rect 2829 36420 2885 36422
rect 2909 36420 2965 36422
rect 6096 36474 6152 36476
rect 6176 36474 6232 36476
rect 6256 36474 6312 36476
rect 6336 36474 6392 36476
rect 6096 36422 6142 36474
rect 6142 36422 6152 36474
rect 6176 36422 6206 36474
rect 6206 36422 6218 36474
rect 6218 36422 6232 36474
rect 6256 36422 6270 36474
rect 6270 36422 6282 36474
rect 6282 36422 6312 36474
rect 6336 36422 6346 36474
rect 6346 36422 6392 36474
rect 6096 36420 6152 36422
rect 6176 36420 6232 36422
rect 6256 36420 6312 36422
rect 6336 36420 6392 36422
rect 9523 36474 9579 36476
rect 9603 36474 9659 36476
rect 9683 36474 9739 36476
rect 9763 36474 9819 36476
rect 9523 36422 9569 36474
rect 9569 36422 9579 36474
rect 9603 36422 9633 36474
rect 9633 36422 9645 36474
rect 9645 36422 9659 36474
rect 9683 36422 9697 36474
rect 9697 36422 9709 36474
rect 9709 36422 9739 36474
rect 9763 36422 9773 36474
rect 9773 36422 9819 36474
rect 9523 36420 9579 36422
rect 9603 36420 9659 36422
rect 9683 36420 9739 36422
rect 9763 36420 9819 36422
rect 12950 36474 13006 36476
rect 13030 36474 13086 36476
rect 13110 36474 13166 36476
rect 13190 36474 13246 36476
rect 12950 36422 12996 36474
rect 12996 36422 13006 36474
rect 13030 36422 13060 36474
rect 13060 36422 13072 36474
rect 13072 36422 13086 36474
rect 13110 36422 13124 36474
rect 13124 36422 13136 36474
rect 13136 36422 13166 36474
rect 13190 36422 13200 36474
rect 13200 36422 13246 36474
rect 12950 36420 13006 36422
rect 13030 36420 13086 36422
rect 13110 36420 13166 36422
rect 13190 36420 13246 36422
rect 4382 35930 4438 35932
rect 4462 35930 4518 35932
rect 4542 35930 4598 35932
rect 4622 35930 4678 35932
rect 4382 35878 4428 35930
rect 4428 35878 4438 35930
rect 4462 35878 4492 35930
rect 4492 35878 4504 35930
rect 4504 35878 4518 35930
rect 4542 35878 4556 35930
rect 4556 35878 4568 35930
rect 4568 35878 4598 35930
rect 4622 35878 4632 35930
rect 4632 35878 4678 35930
rect 4382 35876 4438 35878
rect 4462 35876 4518 35878
rect 4542 35876 4598 35878
rect 4622 35876 4678 35878
rect 7809 35930 7865 35932
rect 7889 35930 7945 35932
rect 7969 35930 8025 35932
rect 8049 35930 8105 35932
rect 7809 35878 7855 35930
rect 7855 35878 7865 35930
rect 7889 35878 7919 35930
rect 7919 35878 7931 35930
rect 7931 35878 7945 35930
rect 7969 35878 7983 35930
rect 7983 35878 7995 35930
rect 7995 35878 8025 35930
rect 8049 35878 8059 35930
rect 8059 35878 8105 35930
rect 7809 35876 7865 35878
rect 7889 35876 7945 35878
rect 7969 35876 8025 35878
rect 8049 35876 8105 35878
rect 11236 35930 11292 35932
rect 11316 35930 11372 35932
rect 11396 35930 11452 35932
rect 11476 35930 11532 35932
rect 11236 35878 11282 35930
rect 11282 35878 11292 35930
rect 11316 35878 11346 35930
rect 11346 35878 11358 35930
rect 11358 35878 11372 35930
rect 11396 35878 11410 35930
rect 11410 35878 11422 35930
rect 11422 35878 11452 35930
rect 11476 35878 11486 35930
rect 11486 35878 11532 35930
rect 11236 35876 11292 35878
rect 11316 35876 11372 35878
rect 11396 35876 11452 35878
rect 11476 35876 11532 35878
rect 14663 35930 14719 35932
rect 14743 35930 14799 35932
rect 14823 35930 14879 35932
rect 14903 35930 14959 35932
rect 14663 35878 14709 35930
rect 14709 35878 14719 35930
rect 14743 35878 14773 35930
rect 14773 35878 14785 35930
rect 14785 35878 14799 35930
rect 14823 35878 14837 35930
rect 14837 35878 14849 35930
rect 14849 35878 14879 35930
rect 14903 35878 14913 35930
rect 14913 35878 14959 35930
rect 14663 35876 14719 35878
rect 14743 35876 14799 35878
rect 14823 35876 14879 35878
rect 14903 35876 14959 35878
rect 14462 35672 14518 35728
rect 2669 35386 2725 35388
rect 2749 35386 2805 35388
rect 2829 35386 2885 35388
rect 2909 35386 2965 35388
rect 2669 35334 2715 35386
rect 2715 35334 2725 35386
rect 2749 35334 2779 35386
rect 2779 35334 2791 35386
rect 2791 35334 2805 35386
rect 2829 35334 2843 35386
rect 2843 35334 2855 35386
rect 2855 35334 2885 35386
rect 2909 35334 2919 35386
rect 2919 35334 2965 35386
rect 2669 35332 2725 35334
rect 2749 35332 2805 35334
rect 2829 35332 2885 35334
rect 2909 35332 2965 35334
rect 6096 35386 6152 35388
rect 6176 35386 6232 35388
rect 6256 35386 6312 35388
rect 6336 35386 6392 35388
rect 6096 35334 6142 35386
rect 6142 35334 6152 35386
rect 6176 35334 6206 35386
rect 6206 35334 6218 35386
rect 6218 35334 6232 35386
rect 6256 35334 6270 35386
rect 6270 35334 6282 35386
rect 6282 35334 6312 35386
rect 6336 35334 6346 35386
rect 6346 35334 6392 35386
rect 6096 35332 6152 35334
rect 6176 35332 6232 35334
rect 6256 35332 6312 35334
rect 6336 35332 6392 35334
rect 9523 35386 9579 35388
rect 9603 35386 9659 35388
rect 9683 35386 9739 35388
rect 9763 35386 9819 35388
rect 9523 35334 9569 35386
rect 9569 35334 9579 35386
rect 9603 35334 9633 35386
rect 9633 35334 9645 35386
rect 9645 35334 9659 35386
rect 9683 35334 9697 35386
rect 9697 35334 9709 35386
rect 9709 35334 9739 35386
rect 9763 35334 9773 35386
rect 9773 35334 9819 35386
rect 9523 35332 9579 35334
rect 9603 35332 9659 35334
rect 9683 35332 9739 35334
rect 9763 35332 9819 35334
rect 12950 35386 13006 35388
rect 13030 35386 13086 35388
rect 13110 35386 13166 35388
rect 13190 35386 13246 35388
rect 12950 35334 12996 35386
rect 12996 35334 13006 35386
rect 13030 35334 13060 35386
rect 13060 35334 13072 35386
rect 13072 35334 13086 35386
rect 13110 35334 13124 35386
rect 13124 35334 13136 35386
rect 13136 35334 13166 35386
rect 13190 35334 13200 35386
rect 13200 35334 13246 35386
rect 12950 35332 13006 35334
rect 13030 35332 13086 35334
rect 13110 35332 13166 35334
rect 13190 35332 13246 35334
rect 4382 34842 4438 34844
rect 4462 34842 4518 34844
rect 4542 34842 4598 34844
rect 4622 34842 4678 34844
rect 4382 34790 4428 34842
rect 4428 34790 4438 34842
rect 4462 34790 4492 34842
rect 4492 34790 4504 34842
rect 4504 34790 4518 34842
rect 4542 34790 4556 34842
rect 4556 34790 4568 34842
rect 4568 34790 4598 34842
rect 4622 34790 4632 34842
rect 4632 34790 4678 34842
rect 4382 34788 4438 34790
rect 4462 34788 4518 34790
rect 4542 34788 4598 34790
rect 4622 34788 4678 34790
rect 7809 34842 7865 34844
rect 7889 34842 7945 34844
rect 7969 34842 8025 34844
rect 8049 34842 8105 34844
rect 7809 34790 7855 34842
rect 7855 34790 7865 34842
rect 7889 34790 7919 34842
rect 7919 34790 7931 34842
rect 7931 34790 7945 34842
rect 7969 34790 7983 34842
rect 7983 34790 7995 34842
rect 7995 34790 8025 34842
rect 8049 34790 8059 34842
rect 8059 34790 8105 34842
rect 7809 34788 7865 34790
rect 7889 34788 7945 34790
rect 7969 34788 8025 34790
rect 8049 34788 8105 34790
rect 11236 34842 11292 34844
rect 11316 34842 11372 34844
rect 11396 34842 11452 34844
rect 11476 34842 11532 34844
rect 11236 34790 11282 34842
rect 11282 34790 11292 34842
rect 11316 34790 11346 34842
rect 11346 34790 11358 34842
rect 11358 34790 11372 34842
rect 11396 34790 11410 34842
rect 11410 34790 11422 34842
rect 11422 34790 11452 34842
rect 11476 34790 11486 34842
rect 11486 34790 11532 34842
rect 11236 34788 11292 34790
rect 11316 34788 11372 34790
rect 11396 34788 11452 34790
rect 11476 34788 11532 34790
rect 14663 34842 14719 34844
rect 14743 34842 14799 34844
rect 14823 34842 14879 34844
rect 14903 34842 14959 34844
rect 14663 34790 14709 34842
rect 14709 34790 14719 34842
rect 14743 34790 14773 34842
rect 14773 34790 14785 34842
rect 14785 34790 14799 34842
rect 14823 34790 14837 34842
rect 14837 34790 14849 34842
rect 14849 34790 14879 34842
rect 14903 34790 14913 34842
rect 14913 34790 14959 34842
rect 14663 34788 14719 34790
rect 14743 34788 14799 34790
rect 14823 34788 14879 34790
rect 14903 34788 14959 34790
rect 2669 34298 2725 34300
rect 2749 34298 2805 34300
rect 2829 34298 2885 34300
rect 2909 34298 2965 34300
rect 2669 34246 2715 34298
rect 2715 34246 2725 34298
rect 2749 34246 2779 34298
rect 2779 34246 2791 34298
rect 2791 34246 2805 34298
rect 2829 34246 2843 34298
rect 2843 34246 2855 34298
rect 2855 34246 2885 34298
rect 2909 34246 2919 34298
rect 2919 34246 2965 34298
rect 2669 34244 2725 34246
rect 2749 34244 2805 34246
rect 2829 34244 2885 34246
rect 2909 34244 2965 34246
rect 6096 34298 6152 34300
rect 6176 34298 6232 34300
rect 6256 34298 6312 34300
rect 6336 34298 6392 34300
rect 6096 34246 6142 34298
rect 6142 34246 6152 34298
rect 6176 34246 6206 34298
rect 6206 34246 6218 34298
rect 6218 34246 6232 34298
rect 6256 34246 6270 34298
rect 6270 34246 6282 34298
rect 6282 34246 6312 34298
rect 6336 34246 6346 34298
rect 6346 34246 6392 34298
rect 6096 34244 6152 34246
rect 6176 34244 6232 34246
rect 6256 34244 6312 34246
rect 6336 34244 6392 34246
rect 9523 34298 9579 34300
rect 9603 34298 9659 34300
rect 9683 34298 9739 34300
rect 9763 34298 9819 34300
rect 9523 34246 9569 34298
rect 9569 34246 9579 34298
rect 9603 34246 9633 34298
rect 9633 34246 9645 34298
rect 9645 34246 9659 34298
rect 9683 34246 9697 34298
rect 9697 34246 9709 34298
rect 9709 34246 9739 34298
rect 9763 34246 9773 34298
rect 9773 34246 9819 34298
rect 9523 34244 9579 34246
rect 9603 34244 9659 34246
rect 9683 34244 9739 34246
rect 9763 34244 9819 34246
rect 12950 34298 13006 34300
rect 13030 34298 13086 34300
rect 13110 34298 13166 34300
rect 13190 34298 13246 34300
rect 12950 34246 12996 34298
rect 12996 34246 13006 34298
rect 13030 34246 13060 34298
rect 13060 34246 13072 34298
rect 13072 34246 13086 34298
rect 13110 34246 13124 34298
rect 13124 34246 13136 34298
rect 13136 34246 13166 34298
rect 13190 34246 13200 34298
rect 13200 34246 13246 34298
rect 12950 34244 13006 34246
rect 13030 34244 13086 34246
rect 13110 34244 13166 34246
rect 13190 34244 13246 34246
rect 4382 33754 4438 33756
rect 4462 33754 4518 33756
rect 4542 33754 4598 33756
rect 4622 33754 4678 33756
rect 4382 33702 4428 33754
rect 4428 33702 4438 33754
rect 4462 33702 4492 33754
rect 4492 33702 4504 33754
rect 4504 33702 4518 33754
rect 4542 33702 4556 33754
rect 4556 33702 4568 33754
rect 4568 33702 4598 33754
rect 4622 33702 4632 33754
rect 4632 33702 4678 33754
rect 4382 33700 4438 33702
rect 4462 33700 4518 33702
rect 4542 33700 4598 33702
rect 4622 33700 4678 33702
rect 7809 33754 7865 33756
rect 7889 33754 7945 33756
rect 7969 33754 8025 33756
rect 8049 33754 8105 33756
rect 7809 33702 7855 33754
rect 7855 33702 7865 33754
rect 7889 33702 7919 33754
rect 7919 33702 7931 33754
rect 7931 33702 7945 33754
rect 7969 33702 7983 33754
rect 7983 33702 7995 33754
rect 7995 33702 8025 33754
rect 8049 33702 8059 33754
rect 8059 33702 8105 33754
rect 7809 33700 7865 33702
rect 7889 33700 7945 33702
rect 7969 33700 8025 33702
rect 8049 33700 8105 33702
rect 11236 33754 11292 33756
rect 11316 33754 11372 33756
rect 11396 33754 11452 33756
rect 11476 33754 11532 33756
rect 11236 33702 11282 33754
rect 11282 33702 11292 33754
rect 11316 33702 11346 33754
rect 11346 33702 11358 33754
rect 11358 33702 11372 33754
rect 11396 33702 11410 33754
rect 11410 33702 11422 33754
rect 11422 33702 11452 33754
rect 11476 33702 11486 33754
rect 11486 33702 11532 33754
rect 11236 33700 11292 33702
rect 11316 33700 11372 33702
rect 11396 33700 11452 33702
rect 11476 33700 11532 33702
rect 14663 33754 14719 33756
rect 14743 33754 14799 33756
rect 14823 33754 14879 33756
rect 14903 33754 14959 33756
rect 14663 33702 14709 33754
rect 14709 33702 14719 33754
rect 14743 33702 14773 33754
rect 14773 33702 14785 33754
rect 14785 33702 14799 33754
rect 14823 33702 14837 33754
rect 14837 33702 14849 33754
rect 14849 33702 14879 33754
rect 14903 33702 14913 33754
rect 14913 33702 14959 33754
rect 14663 33700 14719 33702
rect 14743 33700 14799 33702
rect 14823 33700 14879 33702
rect 14903 33700 14959 33702
rect 2669 33210 2725 33212
rect 2749 33210 2805 33212
rect 2829 33210 2885 33212
rect 2909 33210 2965 33212
rect 2669 33158 2715 33210
rect 2715 33158 2725 33210
rect 2749 33158 2779 33210
rect 2779 33158 2791 33210
rect 2791 33158 2805 33210
rect 2829 33158 2843 33210
rect 2843 33158 2855 33210
rect 2855 33158 2885 33210
rect 2909 33158 2919 33210
rect 2919 33158 2965 33210
rect 2669 33156 2725 33158
rect 2749 33156 2805 33158
rect 2829 33156 2885 33158
rect 2909 33156 2965 33158
rect 6096 33210 6152 33212
rect 6176 33210 6232 33212
rect 6256 33210 6312 33212
rect 6336 33210 6392 33212
rect 6096 33158 6142 33210
rect 6142 33158 6152 33210
rect 6176 33158 6206 33210
rect 6206 33158 6218 33210
rect 6218 33158 6232 33210
rect 6256 33158 6270 33210
rect 6270 33158 6282 33210
rect 6282 33158 6312 33210
rect 6336 33158 6346 33210
rect 6346 33158 6392 33210
rect 6096 33156 6152 33158
rect 6176 33156 6232 33158
rect 6256 33156 6312 33158
rect 6336 33156 6392 33158
rect 9523 33210 9579 33212
rect 9603 33210 9659 33212
rect 9683 33210 9739 33212
rect 9763 33210 9819 33212
rect 9523 33158 9569 33210
rect 9569 33158 9579 33210
rect 9603 33158 9633 33210
rect 9633 33158 9645 33210
rect 9645 33158 9659 33210
rect 9683 33158 9697 33210
rect 9697 33158 9709 33210
rect 9709 33158 9739 33210
rect 9763 33158 9773 33210
rect 9773 33158 9819 33210
rect 9523 33156 9579 33158
rect 9603 33156 9659 33158
rect 9683 33156 9739 33158
rect 9763 33156 9819 33158
rect 12950 33210 13006 33212
rect 13030 33210 13086 33212
rect 13110 33210 13166 33212
rect 13190 33210 13246 33212
rect 12950 33158 12996 33210
rect 12996 33158 13006 33210
rect 13030 33158 13060 33210
rect 13060 33158 13072 33210
rect 13072 33158 13086 33210
rect 13110 33158 13124 33210
rect 13124 33158 13136 33210
rect 13136 33158 13166 33210
rect 13190 33158 13200 33210
rect 13200 33158 13246 33210
rect 12950 33156 13006 33158
rect 13030 33156 13086 33158
rect 13110 33156 13166 33158
rect 13190 33156 13246 33158
rect 4382 32666 4438 32668
rect 4462 32666 4518 32668
rect 4542 32666 4598 32668
rect 4622 32666 4678 32668
rect 4382 32614 4428 32666
rect 4428 32614 4438 32666
rect 4462 32614 4492 32666
rect 4492 32614 4504 32666
rect 4504 32614 4518 32666
rect 4542 32614 4556 32666
rect 4556 32614 4568 32666
rect 4568 32614 4598 32666
rect 4622 32614 4632 32666
rect 4632 32614 4678 32666
rect 4382 32612 4438 32614
rect 4462 32612 4518 32614
rect 4542 32612 4598 32614
rect 4622 32612 4678 32614
rect 7809 32666 7865 32668
rect 7889 32666 7945 32668
rect 7969 32666 8025 32668
rect 8049 32666 8105 32668
rect 7809 32614 7855 32666
rect 7855 32614 7865 32666
rect 7889 32614 7919 32666
rect 7919 32614 7931 32666
rect 7931 32614 7945 32666
rect 7969 32614 7983 32666
rect 7983 32614 7995 32666
rect 7995 32614 8025 32666
rect 8049 32614 8059 32666
rect 8059 32614 8105 32666
rect 7809 32612 7865 32614
rect 7889 32612 7945 32614
rect 7969 32612 8025 32614
rect 8049 32612 8105 32614
rect 11236 32666 11292 32668
rect 11316 32666 11372 32668
rect 11396 32666 11452 32668
rect 11476 32666 11532 32668
rect 11236 32614 11282 32666
rect 11282 32614 11292 32666
rect 11316 32614 11346 32666
rect 11346 32614 11358 32666
rect 11358 32614 11372 32666
rect 11396 32614 11410 32666
rect 11410 32614 11422 32666
rect 11422 32614 11452 32666
rect 11476 32614 11486 32666
rect 11486 32614 11532 32666
rect 11236 32612 11292 32614
rect 11316 32612 11372 32614
rect 11396 32612 11452 32614
rect 11476 32612 11532 32614
rect 14663 32666 14719 32668
rect 14743 32666 14799 32668
rect 14823 32666 14879 32668
rect 14903 32666 14959 32668
rect 14663 32614 14709 32666
rect 14709 32614 14719 32666
rect 14743 32614 14773 32666
rect 14773 32614 14785 32666
rect 14785 32614 14799 32666
rect 14823 32614 14837 32666
rect 14837 32614 14849 32666
rect 14849 32614 14879 32666
rect 14903 32614 14913 32666
rect 14913 32614 14959 32666
rect 14663 32612 14719 32614
rect 14743 32612 14799 32614
rect 14823 32612 14879 32614
rect 14903 32612 14959 32614
rect 2669 32122 2725 32124
rect 2749 32122 2805 32124
rect 2829 32122 2885 32124
rect 2909 32122 2965 32124
rect 2669 32070 2715 32122
rect 2715 32070 2725 32122
rect 2749 32070 2779 32122
rect 2779 32070 2791 32122
rect 2791 32070 2805 32122
rect 2829 32070 2843 32122
rect 2843 32070 2855 32122
rect 2855 32070 2885 32122
rect 2909 32070 2919 32122
rect 2919 32070 2965 32122
rect 2669 32068 2725 32070
rect 2749 32068 2805 32070
rect 2829 32068 2885 32070
rect 2909 32068 2965 32070
rect 6096 32122 6152 32124
rect 6176 32122 6232 32124
rect 6256 32122 6312 32124
rect 6336 32122 6392 32124
rect 6096 32070 6142 32122
rect 6142 32070 6152 32122
rect 6176 32070 6206 32122
rect 6206 32070 6218 32122
rect 6218 32070 6232 32122
rect 6256 32070 6270 32122
rect 6270 32070 6282 32122
rect 6282 32070 6312 32122
rect 6336 32070 6346 32122
rect 6346 32070 6392 32122
rect 6096 32068 6152 32070
rect 6176 32068 6232 32070
rect 6256 32068 6312 32070
rect 6336 32068 6392 32070
rect 9523 32122 9579 32124
rect 9603 32122 9659 32124
rect 9683 32122 9739 32124
rect 9763 32122 9819 32124
rect 9523 32070 9569 32122
rect 9569 32070 9579 32122
rect 9603 32070 9633 32122
rect 9633 32070 9645 32122
rect 9645 32070 9659 32122
rect 9683 32070 9697 32122
rect 9697 32070 9709 32122
rect 9709 32070 9739 32122
rect 9763 32070 9773 32122
rect 9773 32070 9819 32122
rect 9523 32068 9579 32070
rect 9603 32068 9659 32070
rect 9683 32068 9739 32070
rect 9763 32068 9819 32070
rect 12950 32122 13006 32124
rect 13030 32122 13086 32124
rect 13110 32122 13166 32124
rect 13190 32122 13246 32124
rect 12950 32070 12996 32122
rect 12996 32070 13006 32122
rect 13030 32070 13060 32122
rect 13060 32070 13072 32122
rect 13072 32070 13086 32122
rect 13110 32070 13124 32122
rect 13124 32070 13136 32122
rect 13136 32070 13166 32122
rect 13190 32070 13200 32122
rect 13200 32070 13246 32122
rect 12950 32068 13006 32070
rect 13030 32068 13086 32070
rect 13110 32068 13166 32070
rect 13190 32068 13246 32070
rect 4382 31578 4438 31580
rect 4462 31578 4518 31580
rect 4542 31578 4598 31580
rect 4622 31578 4678 31580
rect 4382 31526 4428 31578
rect 4428 31526 4438 31578
rect 4462 31526 4492 31578
rect 4492 31526 4504 31578
rect 4504 31526 4518 31578
rect 4542 31526 4556 31578
rect 4556 31526 4568 31578
rect 4568 31526 4598 31578
rect 4622 31526 4632 31578
rect 4632 31526 4678 31578
rect 4382 31524 4438 31526
rect 4462 31524 4518 31526
rect 4542 31524 4598 31526
rect 4622 31524 4678 31526
rect 7809 31578 7865 31580
rect 7889 31578 7945 31580
rect 7969 31578 8025 31580
rect 8049 31578 8105 31580
rect 7809 31526 7855 31578
rect 7855 31526 7865 31578
rect 7889 31526 7919 31578
rect 7919 31526 7931 31578
rect 7931 31526 7945 31578
rect 7969 31526 7983 31578
rect 7983 31526 7995 31578
rect 7995 31526 8025 31578
rect 8049 31526 8059 31578
rect 8059 31526 8105 31578
rect 7809 31524 7865 31526
rect 7889 31524 7945 31526
rect 7969 31524 8025 31526
rect 8049 31524 8105 31526
rect 11236 31578 11292 31580
rect 11316 31578 11372 31580
rect 11396 31578 11452 31580
rect 11476 31578 11532 31580
rect 11236 31526 11282 31578
rect 11282 31526 11292 31578
rect 11316 31526 11346 31578
rect 11346 31526 11358 31578
rect 11358 31526 11372 31578
rect 11396 31526 11410 31578
rect 11410 31526 11422 31578
rect 11422 31526 11452 31578
rect 11476 31526 11486 31578
rect 11486 31526 11532 31578
rect 11236 31524 11292 31526
rect 11316 31524 11372 31526
rect 11396 31524 11452 31526
rect 11476 31524 11532 31526
rect 14663 31578 14719 31580
rect 14743 31578 14799 31580
rect 14823 31578 14879 31580
rect 14903 31578 14959 31580
rect 14663 31526 14709 31578
rect 14709 31526 14719 31578
rect 14743 31526 14773 31578
rect 14773 31526 14785 31578
rect 14785 31526 14799 31578
rect 14823 31526 14837 31578
rect 14837 31526 14849 31578
rect 14849 31526 14879 31578
rect 14903 31526 14913 31578
rect 14913 31526 14959 31578
rect 14663 31524 14719 31526
rect 14743 31524 14799 31526
rect 14823 31524 14879 31526
rect 14903 31524 14959 31526
rect 2669 31034 2725 31036
rect 2749 31034 2805 31036
rect 2829 31034 2885 31036
rect 2909 31034 2965 31036
rect 2669 30982 2715 31034
rect 2715 30982 2725 31034
rect 2749 30982 2779 31034
rect 2779 30982 2791 31034
rect 2791 30982 2805 31034
rect 2829 30982 2843 31034
rect 2843 30982 2855 31034
rect 2855 30982 2885 31034
rect 2909 30982 2919 31034
rect 2919 30982 2965 31034
rect 2669 30980 2725 30982
rect 2749 30980 2805 30982
rect 2829 30980 2885 30982
rect 2909 30980 2965 30982
rect 6096 31034 6152 31036
rect 6176 31034 6232 31036
rect 6256 31034 6312 31036
rect 6336 31034 6392 31036
rect 6096 30982 6142 31034
rect 6142 30982 6152 31034
rect 6176 30982 6206 31034
rect 6206 30982 6218 31034
rect 6218 30982 6232 31034
rect 6256 30982 6270 31034
rect 6270 30982 6282 31034
rect 6282 30982 6312 31034
rect 6336 30982 6346 31034
rect 6346 30982 6392 31034
rect 6096 30980 6152 30982
rect 6176 30980 6232 30982
rect 6256 30980 6312 30982
rect 6336 30980 6392 30982
rect 9523 31034 9579 31036
rect 9603 31034 9659 31036
rect 9683 31034 9739 31036
rect 9763 31034 9819 31036
rect 9523 30982 9569 31034
rect 9569 30982 9579 31034
rect 9603 30982 9633 31034
rect 9633 30982 9645 31034
rect 9645 30982 9659 31034
rect 9683 30982 9697 31034
rect 9697 30982 9709 31034
rect 9709 30982 9739 31034
rect 9763 30982 9773 31034
rect 9773 30982 9819 31034
rect 9523 30980 9579 30982
rect 9603 30980 9659 30982
rect 9683 30980 9739 30982
rect 9763 30980 9819 30982
rect 12950 31034 13006 31036
rect 13030 31034 13086 31036
rect 13110 31034 13166 31036
rect 13190 31034 13246 31036
rect 12950 30982 12996 31034
rect 12996 30982 13006 31034
rect 13030 30982 13060 31034
rect 13060 30982 13072 31034
rect 13072 30982 13086 31034
rect 13110 30982 13124 31034
rect 13124 30982 13136 31034
rect 13136 30982 13166 31034
rect 13190 30982 13200 31034
rect 13200 30982 13246 31034
rect 12950 30980 13006 30982
rect 13030 30980 13086 30982
rect 13110 30980 13166 30982
rect 13190 30980 13246 30982
rect 4382 30490 4438 30492
rect 4462 30490 4518 30492
rect 4542 30490 4598 30492
rect 4622 30490 4678 30492
rect 4382 30438 4428 30490
rect 4428 30438 4438 30490
rect 4462 30438 4492 30490
rect 4492 30438 4504 30490
rect 4504 30438 4518 30490
rect 4542 30438 4556 30490
rect 4556 30438 4568 30490
rect 4568 30438 4598 30490
rect 4622 30438 4632 30490
rect 4632 30438 4678 30490
rect 4382 30436 4438 30438
rect 4462 30436 4518 30438
rect 4542 30436 4598 30438
rect 4622 30436 4678 30438
rect 7809 30490 7865 30492
rect 7889 30490 7945 30492
rect 7969 30490 8025 30492
rect 8049 30490 8105 30492
rect 7809 30438 7855 30490
rect 7855 30438 7865 30490
rect 7889 30438 7919 30490
rect 7919 30438 7931 30490
rect 7931 30438 7945 30490
rect 7969 30438 7983 30490
rect 7983 30438 7995 30490
rect 7995 30438 8025 30490
rect 8049 30438 8059 30490
rect 8059 30438 8105 30490
rect 7809 30436 7865 30438
rect 7889 30436 7945 30438
rect 7969 30436 8025 30438
rect 8049 30436 8105 30438
rect 11236 30490 11292 30492
rect 11316 30490 11372 30492
rect 11396 30490 11452 30492
rect 11476 30490 11532 30492
rect 11236 30438 11282 30490
rect 11282 30438 11292 30490
rect 11316 30438 11346 30490
rect 11346 30438 11358 30490
rect 11358 30438 11372 30490
rect 11396 30438 11410 30490
rect 11410 30438 11422 30490
rect 11422 30438 11452 30490
rect 11476 30438 11486 30490
rect 11486 30438 11532 30490
rect 11236 30436 11292 30438
rect 11316 30436 11372 30438
rect 11396 30436 11452 30438
rect 11476 30436 11532 30438
rect 14663 30490 14719 30492
rect 14743 30490 14799 30492
rect 14823 30490 14879 30492
rect 14903 30490 14959 30492
rect 14663 30438 14709 30490
rect 14709 30438 14719 30490
rect 14743 30438 14773 30490
rect 14773 30438 14785 30490
rect 14785 30438 14799 30490
rect 14823 30438 14837 30490
rect 14837 30438 14849 30490
rect 14849 30438 14879 30490
rect 14903 30438 14913 30490
rect 14913 30438 14959 30490
rect 14663 30436 14719 30438
rect 14743 30436 14799 30438
rect 14823 30436 14879 30438
rect 14903 30436 14959 30438
rect 2669 29946 2725 29948
rect 2749 29946 2805 29948
rect 2829 29946 2885 29948
rect 2909 29946 2965 29948
rect 2669 29894 2715 29946
rect 2715 29894 2725 29946
rect 2749 29894 2779 29946
rect 2779 29894 2791 29946
rect 2791 29894 2805 29946
rect 2829 29894 2843 29946
rect 2843 29894 2855 29946
rect 2855 29894 2885 29946
rect 2909 29894 2919 29946
rect 2919 29894 2965 29946
rect 2669 29892 2725 29894
rect 2749 29892 2805 29894
rect 2829 29892 2885 29894
rect 2909 29892 2965 29894
rect 6096 29946 6152 29948
rect 6176 29946 6232 29948
rect 6256 29946 6312 29948
rect 6336 29946 6392 29948
rect 6096 29894 6142 29946
rect 6142 29894 6152 29946
rect 6176 29894 6206 29946
rect 6206 29894 6218 29946
rect 6218 29894 6232 29946
rect 6256 29894 6270 29946
rect 6270 29894 6282 29946
rect 6282 29894 6312 29946
rect 6336 29894 6346 29946
rect 6346 29894 6392 29946
rect 6096 29892 6152 29894
rect 6176 29892 6232 29894
rect 6256 29892 6312 29894
rect 6336 29892 6392 29894
rect 9523 29946 9579 29948
rect 9603 29946 9659 29948
rect 9683 29946 9739 29948
rect 9763 29946 9819 29948
rect 9523 29894 9569 29946
rect 9569 29894 9579 29946
rect 9603 29894 9633 29946
rect 9633 29894 9645 29946
rect 9645 29894 9659 29946
rect 9683 29894 9697 29946
rect 9697 29894 9709 29946
rect 9709 29894 9739 29946
rect 9763 29894 9773 29946
rect 9773 29894 9819 29946
rect 9523 29892 9579 29894
rect 9603 29892 9659 29894
rect 9683 29892 9739 29894
rect 9763 29892 9819 29894
rect 12950 29946 13006 29948
rect 13030 29946 13086 29948
rect 13110 29946 13166 29948
rect 13190 29946 13246 29948
rect 12950 29894 12996 29946
rect 12996 29894 13006 29946
rect 13030 29894 13060 29946
rect 13060 29894 13072 29946
rect 13072 29894 13086 29946
rect 13110 29894 13124 29946
rect 13124 29894 13136 29946
rect 13136 29894 13166 29946
rect 13190 29894 13200 29946
rect 13200 29894 13246 29946
rect 12950 29892 13006 29894
rect 13030 29892 13086 29894
rect 13110 29892 13166 29894
rect 13190 29892 13246 29894
rect 4382 29402 4438 29404
rect 4462 29402 4518 29404
rect 4542 29402 4598 29404
rect 4622 29402 4678 29404
rect 4382 29350 4428 29402
rect 4428 29350 4438 29402
rect 4462 29350 4492 29402
rect 4492 29350 4504 29402
rect 4504 29350 4518 29402
rect 4542 29350 4556 29402
rect 4556 29350 4568 29402
rect 4568 29350 4598 29402
rect 4622 29350 4632 29402
rect 4632 29350 4678 29402
rect 4382 29348 4438 29350
rect 4462 29348 4518 29350
rect 4542 29348 4598 29350
rect 4622 29348 4678 29350
rect 7809 29402 7865 29404
rect 7889 29402 7945 29404
rect 7969 29402 8025 29404
rect 8049 29402 8105 29404
rect 7809 29350 7855 29402
rect 7855 29350 7865 29402
rect 7889 29350 7919 29402
rect 7919 29350 7931 29402
rect 7931 29350 7945 29402
rect 7969 29350 7983 29402
rect 7983 29350 7995 29402
rect 7995 29350 8025 29402
rect 8049 29350 8059 29402
rect 8059 29350 8105 29402
rect 7809 29348 7865 29350
rect 7889 29348 7945 29350
rect 7969 29348 8025 29350
rect 8049 29348 8105 29350
rect 11236 29402 11292 29404
rect 11316 29402 11372 29404
rect 11396 29402 11452 29404
rect 11476 29402 11532 29404
rect 11236 29350 11282 29402
rect 11282 29350 11292 29402
rect 11316 29350 11346 29402
rect 11346 29350 11358 29402
rect 11358 29350 11372 29402
rect 11396 29350 11410 29402
rect 11410 29350 11422 29402
rect 11422 29350 11452 29402
rect 11476 29350 11486 29402
rect 11486 29350 11532 29402
rect 11236 29348 11292 29350
rect 11316 29348 11372 29350
rect 11396 29348 11452 29350
rect 11476 29348 11532 29350
rect 14663 29402 14719 29404
rect 14743 29402 14799 29404
rect 14823 29402 14879 29404
rect 14903 29402 14959 29404
rect 14663 29350 14709 29402
rect 14709 29350 14719 29402
rect 14743 29350 14773 29402
rect 14773 29350 14785 29402
rect 14785 29350 14799 29402
rect 14823 29350 14837 29402
rect 14837 29350 14849 29402
rect 14849 29350 14879 29402
rect 14903 29350 14913 29402
rect 14913 29350 14959 29402
rect 14663 29348 14719 29350
rect 14743 29348 14799 29350
rect 14823 29348 14879 29350
rect 14903 29348 14959 29350
rect 2669 28858 2725 28860
rect 2749 28858 2805 28860
rect 2829 28858 2885 28860
rect 2909 28858 2965 28860
rect 2669 28806 2715 28858
rect 2715 28806 2725 28858
rect 2749 28806 2779 28858
rect 2779 28806 2791 28858
rect 2791 28806 2805 28858
rect 2829 28806 2843 28858
rect 2843 28806 2855 28858
rect 2855 28806 2885 28858
rect 2909 28806 2919 28858
rect 2919 28806 2965 28858
rect 2669 28804 2725 28806
rect 2749 28804 2805 28806
rect 2829 28804 2885 28806
rect 2909 28804 2965 28806
rect 6096 28858 6152 28860
rect 6176 28858 6232 28860
rect 6256 28858 6312 28860
rect 6336 28858 6392 28860
rect 6096 28806 6142 28858
rect 6142 28806 6152 28858
rect 6176 28806 6206 28858
rect 6206 28806 6218 28858
rect 6218 28806 6232 28858
rect 6256 28806 6270 28858
rect 6270 28806 6282 28858
rect 6282 28806 6312 28858
rect 6336 28806 6346 28858
rect 6346 28806 6392 28858
rect 6096 28804 6152 28806
rect 6176 28804 6232 28806
rect 6256 28804 6312 28806
rect 6336 28804 6392 28806
rect 9523 28858 9579 28860
rect 9603 28858 9659 28860
rect 9683 28858 9739 28860
rect 9763 28858 9819 28860
rect 9523 28806 9569 28858
rect 9569 28806 9579 28858
rect 9603 28806 9633 28858
rect 9633 28806 9645 28858
rect 9645 28806 9659 28858
rect 9683 28806 9697 28858
rect 9697 28806 9709 28858
rect 9709 28806 9739 28858
rect 9763 28806 9773 28858
rect 9773 28806 9819 28858
rect 9523 28804 9579 28806
rect 9603 28804 9659 28806
rect 9683 28804 9739 28806
rect 9763 28804 9819 28806
rect 12950 28858 13006 28860
rect 13030 28858 13086 28860
rect 13110 28858 13166 28860
rect 13190 28858 13246 28860
rect 12950 28806 12996 28858
rect 12996 28806 13006 28858
rect 13030 28806 13060 28858
rect 13060 28806 13072 28858
rect 13072 28806 13086 28858
rect 13110 28806 13124 28858
rect 13124 28806 13136 28858
rect 13136 28806 13166 28858
rect 13190 28806 13200 28858
rect 13200 28806 13246 28858
rect 12950 28804 13006 28806
rect 13030 28804 13086 28806
rect 13110 28804 13166 28806
rect 13190 28804 13246 28806
rect 4382 28314 4438 28316
rect 4462 28314 4518 28316
rect 4542 28314 4598 28316
rect 4622 28314 4678 28316
rect 4382 28262 4428 28314
rect 4428 28262 4438 28314
rect 4462 28262 4492 28314
rect 4492 28262 4504 28314
rect 4504 28262 4518 28314
rect 4542 28262 4556 28314
rect 4556 28262 4568 28314
rect 4568 28262 4598 28314
rect 4622 28262 4632 28314
rect 4632 28262 4678 28314
rect 4382 28260 4438 28262
rect 4462 28260 4518 28262
rect 4542 28260 4598 28262
rect 4622 28260 4678 28262
rect 7809 28314 7865 28316
rect 7889 28314 7945 28316
rect 7969 28314 8025 28316
rect 8049 28314 8105 28316
rect 7809 28262 7855 28314
rect 7855 28262 7865 28314
rect 7889 28262 7919 28314
rect 7919 28262 7931 28314
rect 7931 28262 7945 28314
rect 7969 28262 7983 28314
rect 7983 28262 7995 28314
rect 7995 28262 8025 28314
rect 8049 28262 8059 28314
rect 8059 28262 8105 28314
rect 7809 28260 7865 28262
rect 7889 28260 7945 28262
rect 7969 28260 8025 28262
rect 8049 28260 8105 28262
rect 11236 28314 11292 28316
rect 11316 28314 11372 28316
rect 11396 28314 11452 28316
rect 11476 28314 11532 28316
rect 11236 28262 11282 28314
rect 11282 28262 11292 28314
rect 11316 28262 11346 28314
rect 11346 28262 11358 28314
rect 11358 28262 11372 28314
rect 11396 28262 11410 28314
rect 11410 28262 11422 28314
rect 11422 28262 11452 28314
rect 11476 28262 11486 28314
rect 11486 28262 11532 28314
rect 11236 28260 11292 28262
rect 11316 28260 11372 28262
rect 11396 28260 11452 28262
rect 11476 28260 11532 28262
rect 14663 28314 14719 28316
rect 14743 28314 14799 28316
rect 14823 28314 14879 28316
rect 14903 28314 14959 28316
rect 14663 28262 14709 28314
rect 14709 28262 14719 28314
rect 14743 28262 14773 28314
rect 14773 28262 14785 28314
rect 14785 28262 14799 28314
rect 14823 28262 14837 28314
rect 14837 28262 14849 28314
rect 14849 28262 14879 28314
rect 14903 28262 14913 28314
rect 14913 28262 14959 28314
rect 14663 28260 14719 28262
rect 14743 28260 14799 28262
rect 14823 28260 14879 28262
rect 14903 28260 14959 28262
rect 14462 27784 14518 27840
rect 2669 27770 2725 27772
rect 2749 27770 2805 27772
rect 2829 27770 2885 27772
rect 2909 27770 2965 27772
rect 2669 27718 2715 27770
rect 2715 27718 2725 27770
rect 2749 27718 2779 27770
rect 2779 27718 2791 27770
rect 2791 27718 2805 27770
rect 2829 27718 2843 27770
rect 2843 27718 2855 27770
rect 2855 27718 2885 27770
rect 2909 27718 2919 27770
rect 2919 27718 2965 27770
rect 2669 27716 2725 27718
rect 2749 27716 2805 27718
rect 2829 27716 2885 27718
rect 2909 27716 2965 27718
rect 6096 27770 6152 27772
rect 6176 27770 6232 27772
rect 6256 27770 6312 27772
rect 6336 27770 6392 27772
rect 6096 27718 6142 27770
rect 6142 27718 6152 27770
rect 6176 27718 6206 27770
rect 6206 27718 6218 27770
rect 6218 27718 6232 27770
rect 6256 27718 6270 27770
rect 6270 27718 6282 27770
rect 6282 27718 6312 27770
rect 6336 27718 6346 27770
rect 6346 27718 6392 27770
rect 6096 27716 6152 27718
rect 6176 27716 6232 27718
rect 6256 27716 6312 27718
rect 6336 27716 6392 27718
rect 9523 27770 9579 27772
rect 9603 27770 9659 27772
rect 9683 27770 9739 27772
rect 9763 27770 9819 27772
rect 9523 27718 9569 27770
rect 9569 27718 9579 27770
rect 9603 27718 9633 27770
rect 9633 27718 9645 27770
rect 9645 27718 9659 27770
rect 9683 27718 9697 27770
rect 9697 27718 9709 27770
rect 9709 27718 9739 27770
rect 9763 27718 9773 27770
rect 9773 27718 9819 27770
rect 9523 27716 9579 27718
rect 9603 27716 9659 27718
rect 9683 27716 9739 27718
rect 9763 27716 9819 27718
rect 12950 27770 13006 27772
rect 13030 27770 13086 27772
rect 13110 27770 13166 27772
rect 13190 27770 13246 27772
rect 12950 27718 12996 27770
rect 12996 27718 13006 27770
rect 13030 27718 13060 27770
rect 13060 27718 13072 27770
rect 13072 27718 13086 27770
rect 13110 27718 13124 27770
rect 13124 27718 13136 27770
rect 13136 27718 13166 27770
rect 13190 27718 13200 27770
rect 13200 27718 13246 27770
rect 12950 27716 13006 27718
rect 13030 27716 13086 27718
rect 13110 27716 13166 27718
rect 13190 27716 13246 27718
rect 4382 27226 4438 27228
rect 4462 27226 4518 27228
rect 4542 27226 4598 27228
rect 4622 27226 4678 27228
rect 4382 27174 4428 27226
rect 4428 27174 4438 27226
rect 4462 27174 4492 27226
rect 4492 27174 4504 27226
rect 4504 27174 4518 27226
rect 4542 27174 4556 27226
rect 4556 27174 4568 27226
rect 4568 27174 4598 27226
rect 4622 27174 4632 27226
rect 4632 27174 4678 27226
rect 4382 27172 4438 27174
rect 4462 27172 4518 27174
rect 4542 27172 4598 27174
rect 4622 27172 4678 27174
rect 7809 27226 7865 27228
rect 7889 27226 7945 27228
rect 7969 27226 8025 27228
rect 8049 27226 8105 27228
rect 7809 27174 7855 27226
rect 7855 27174 7865 27226
rect 7889 27174 7919 27226
rect 7919 27174 7931 27226
rect 7931 27174 7945 27226
rect 7969 27174 7983 27226
rect 7983 27174 7995 27226
rect 7995 27174 8025 27226
rect 8049 27174 8059 27226
rect 8059 27174 8105 27226
rect 7809 27172 7865 27174
rect 7889 27172 7945 27174
rect 7969 27172 8025 27174
rect 8049 27172 8105 27174
rect 11236 27226 11292 27228
rect 11316 27226 11372 27228
rect 11396 27226 11452 27228
rect 11476 27226 11532 27228
rect 11236 27174 11282 27226
rect 11282 27174 11292 27226
rect 11316 27174 11346 27226
rect 11346 27174 11358 27226
rect 11358 27174 11372 27226
rect 11396 27174 11410 27226
rect 11410 27174 11422 27226
rect 11422 27174 11452 27226
rect 11476 27174 11486 27226
rect 11486 27174 11532 27226
rect 11236 27172 11292 27174
rect 11316 27172 11372 27174
rect 11396 27172 11452 27174
rect 11476 27172 11532 27174
rect 14663 27226 14719 27228
rect 14743 27226 14799 27228
rect 14823 27226 14879 27228
rect 14903 27226 14959 27228
rect 14663 27174 14709 27226
rect 14709 27174 14719 27226
rect 14743 27174 14773 27226
rect 14773 27174 14785 27226
rect 14785 27174 14799 27226
rect 14823 27174 14837 27226
rect 14837 27174 14849 27226
rect 14849 27174 14879 27226
rect 14903 27174 14913 27226
rect 14913 27174 14959 27226
rect 14663 27172 14719 27174
rect 14743 27172 14799 27174
rect 14823 27172 14879 27174
rect 14903 27172 14959 27174
rect 2669 26682 2725 26684
rect 2749 26682 2805 26684
rect 2829 26682 2885 26684
rect 2909 26682 2965 26684
rect 2669 26630 2715 26682
rect 2715 26630 2725 26682
rect 2749 26630 2779 26682
rect 2779 26630 2791 26682
rect 2791 26630 2805 26682
rect 2829 26630 2843 26682
rect 2843 26630 2855 26682
rect 2855 26630 2885 26682
rect 2909 26630 2919 26682
rect 2919 26630 2965 26682
rect 2669 26628 2725 26630
rect 2749 26628 2805 26630
rect 2829 26628 2885 26630
rect 2909 26628 2965 26630
rect 6096 26682 6152 26684
rect 6176 26682 6232 26684
rect 6256 26682 6312 26684
rect 6336 26682 6392 26684
rect 6096 26630 6142 26682
rect 6142 26630 6152 26682
rect 6176 26630 6206 26682
rect 6206 26630 6218 26682
rect 6218 26630 6232 26682
rect 6256 26630 6270 26682
rect 6270 26630 6282 26682
rect 6282 26630 6312 26682
rect 6336 26630 6346 26682
rect 6346 26630 6392 26682
rect 6096 26628 6152 26630
rect 6176 26628 6232 26630
rect 6256 26628 6312 26630
rect 6336 26628 6392 26630
rect 9523 26682 9579 26684
rect 9603 26682 9659 26684
rect 9683 26682 9739 26684
rect 9763 26682 9819 26684
rect 9523 26630 9569 26682
rect 9569 26630 9579 26682
rect 9603 26630 9633 26682
rect 9633 26630 9645 26682
rect 9645 26630 9659 26682
rect 9683 26630 9697 26682
rect 9697 26630 9709 26682
rect 9709 26630 9739 26682
rect 9763 26630 9773 26682
rect 9773 26630 9819 26682
rect 9523 26628 9579 26630
rect 9603 26628 9659 26630
rect 9683 26628 9739 26630
rect 9763 26628 9819 26630
rect 12950 26682 13006 26684
rect 13030 26682 13086 26684
rect 13110 26682 13166 26684
rect 13190 26682 13246 26684
rect 12950 26630 12996 26682
rect 12996 26630 13006 26682
rect 13030 26630 13060 26682
rect 13060 26630 13072 26682
rect 13072 26630 13086 26682
rect 13110 26630 13124 26682
rect 13124 26630 13136 26682
rect 13136 26630 13166 26682
rect 13190 26630 13200 26682
rect 13200 26630 13246 26682
rect 12950 26628 13006 26630
rect 13030 26628 13086 26630
rect 13110 26628 13166 26630
rect 13190 26628 13246 26630
rect 4382 26138 4438 26140
rect 4462 26138 4518 26140
rect 4542 26138 4598 26140
rect 4622 26138 4678 26140
rect 4382 26086 4428 26138
rect 4428 26086 4438 26138
rect 4462 26086 4492 26138
rect 4492 26086 4504 26138
rect 4504 26086 4518 26138
rect 4542 26086 4556 26138
rect 4556 26086 4568 26138
rect 4568 26086 4598 26138
rect 4622 26086 4632 26138
rect 4632 26086 4678 26138
rect 4382 26084 4438 26086
rect 4462 26084 4518 26086
rect 4542 26084 4598 26086
rect 4622 26084 4678 26086
rect 7809 26138 7865 26140
rect 7889 26138 7945 26140
rect 7969 26138 8025 26140
rect 8049 26138 8105 26140
rect 7809 26086 7855 26138
rect 7855 26086 7865 26138
rect 7889 26086 7919 26138
rect 7919 26086 7931 26138
rect 7931 26086 7945 26138
rect 7969 26086 7983 26138
rect 7983 26086 7995 26138
rect 7995 26086 8025 26138
rect 8049 26086 8059 26138
rect 8059 26086 8105 26138
rect 7809 26084 7865 26086
rect 7889 26084 7945 26086
rect 7969 26084 8025 26086
rect 8049 26084 8105 26086
rect 11236 26138 11292 26140
rect 11316 26138 11372 26140
rect 11396 26138 11452 26140
rect 11476 26138 11532 26140
rect 11236 26086 11282 26138
rect 11282 26086 11292 26138
rect 11316 26086 11346 26138
rect 11346 26086 11358 26138
rect 11358 26086 11372 26138
rect 11396 26086 11410 26138
rect 11410 26086 11422 26138
rect 11422 26086 11452 26138
rect 11476 26086 11486 26138
rect 11486 26086 11532 26138
rect 11236 26084 11292 26086
rect 11316 26084 11372 26086
rect 11396 26084 11452 26086
rect 11476 26084 11532 26086
rect 14663 26138 14719 26140
rect 14743 26138 14799 26140
rect 14823 26138 14879 26140
rect 14903 26138 14959 26140
rect 14663 26086 14709 26138
rect 14709 26086 14719 26138
rect 14743 26086 14773 26138
rect 14773 26086 14785 26138
rect 14785 26086 14799 26138
rect 14823 26086 14837 26138
rect 14837 26086 14849 26138
rect 14849 26086 14879 26138
rect 14903 26086 14913 26138
rect 14913 26086 14959 26138
rect 14663 26084 14719 26086
rect 14743 26084 14799 26086
rect 14823 26084 14879 26086
rect 14903 26084 14959 26086
rect 2669 25594 2725 25596
rect 2749 25594 2805 25596
rect 2829 25594 2885 25596
rect 2909 25594 2965 25596
rect 2669 25542 2715 25594
rect 2715 25542 2725 25594
rect 2749 25542 2779 25594
rect 2779 25542 2791 25594
rect 2791 25542 2805 25594
rect 2829 25542 2843 25594
rect 2843 25542 2855 25594
rect 2855 25542 2885 25594
rect 2909 25542 2919 25594
rect 2919 25542 2965 25594
rect 2669 25540 2725 25542
rect 2749 25540 2805 25542
rect 2829 25540 2885 25542
rect 2909 25540 2965 25542
rect 6096 25594 6152 25596
rect 6176 25594 6232 25596
rect 6256 25594 6312 25596
rect 6336 25594 6392 25596
rect 6096 25542 6142 25594
rect 6142 25542 6152 25594
rect 6176 25542 6206 25594
rect 6206 25542 6218 25594
rect 6218 25542 6232 25594
rect 6256 25542 6270 25594
rect 6270 25542 6282 25594
rect 6282 25542 6312 25594
rect 6336 25542 6346 25594
rect 6346 25542 6392 25594
rect 6096 25540 6152 25542
rect 6176 25540 6232 25542
rect 6256 25540 6312 25542
rect 6336 25540 6392 25542
rect 9523 25594 9579 25596
rect 9603 25594 9659 25596
rect 9683 25594 9739 25596
rect 9763 25594 9819 25596
rect 9523 25542 9569 25594
rect 9569 25542 9579 25594
rect 9603 25542 9633 25594
rect 9633 25542 9645 25594
rect 9645 25542 9659 25594
rect 9683 25542 9697 25594
rect 9697 25542 9709 25594
rect 9709 25542 9739 25594
rect 9763 25542 9773 25594
rect 9773 25542 9819 25594
rect 9523 25540 9579 25542
rect 9603 25540 9659 25542
rect 9683 25540 9739 25542
rect 9763 25540 9819 25542
rect 12950 25594 13006 25596
rect 13030 25594 13086 25596
rect 13110 25594 13166 25596
rect 13190 25594 13246 25596
rect 12950 25542 12996 25594
rect 12996 25542 13006 25594
rect 13030 25542 13060 25594
rect 13060 25542 13072 25594
rect 13072 25542 13086 25594
rect 13110 25542 13124 25594
rect 13124 25542 13136 25594
rect 13136 25542 13166 25594
rect 13190 25542 13200 25594
rect 13200 25542 13246 25594
rect 12950 25540 13006 25542
rect 13030 25540 13086 25542
rect 13110 25540 13166 25542
rect 13190 25540 13246 25542
rect 4382 25050 4438 25052
rect 4462 25050 4518 25052
rect 4542 25050 4598 25052
rect 4622 25050 4678 25052
rect 4382 24998 4428 25050
rect 4428 24998 4438 25050
rect 4462 24998 4492 25050
rect 4492 24998 4504 25050
rect 4504 24998 4518 25050
rect 4542 24998 4556 25050
rect 4556 24998 4568 25050
rect 4568 24998 4598 25050
rect 4622 24998 4632 25050
rect 4632 24998 4678 25050
rect 4382 24996 4438 24998
rect 4462 24996 4518 24998
rect 4542 24996 4598 24998
rect 4622 24996 4678 24998
rect 7809 25050 7865 25052
rect 7889 25050 7945 25052
rect 7969 25050 8025 25052
rect 8049 25050 8105 25052
rect 7809 24998 7855 25050
rect 7855 24998 7865 25050
rect 7889 24998 7919 25050
rect 7919 24998 7931 25050
rect 7931 24998 7945 25050
rect 7969 24998 7983 25050
rect 7983 24998 7995 25050
rect 7995 24998 8025 25050
rect 8049 24998 8059 25050
rect 8059 24998 8105 25050
rect 7809 24996 7865 24998
rect 7889 24996 7945 24998
rect 7969 24996 8025 24998
rect 8049 24996 8105 24998
rect 11236 25050 11292 25052
rect 11316 25050 11372 25052
rect 11396 25050 11452 25052
rect 11476 25050 11532 25052
rect 11236 24998 11282 25050
rect 11282 24998 11292 25050
rect 11316 24998 11346 25050
rect 11346 24998 11358 25050
rect 11358 24998 11372 25050
rect 11396 24998 11410 25050
rect 11410 24998 11422 25050
rect 11422 24998 11452 25050
rect 11476 24998 11486 25050
rect 11486 24998 11532 25050
rect 11236 24996 11292 24998
rect 11316 24996 11372 24998
rect 11396 24996 11452 24998
rect 11476 24996 11532 24998
rect 14663 25050 14719 25052
rect 14743 25050 14799 25052
rect 14823 25050 14879 25052
rect 14903 25050 14959 25052
rect 14663 24998 14709 25050
rect 14709 24998 14719 25050
rect 14743 24998 14773 25050
rect 14773 24998 14785 25050
rect 14785 24998 14799 25050
rect 14823 24998 14837 25050
rect 14837 24998 14849 25050
rect 14849 24998 14879 25050
rect 14903 24998 14913 25050
rect 14913 24998 14959 25050
rect 14663 24996 14719 24998
rect 14743 24996 14799 24998
rect 14823 24996 14879 24998
rect 14903 24996 14959 24998
rect 2669 24506 2725 24508
rect 2749 24506 2805 24508
rect 2829 24506 2885 24508
rect 2909 24506 2965 24508
rect 2669 24454 2715 24506
rect 2715 24454 2725 24506
rect 2749 24454 2779 24506
rect 2779 24454 2791 24506
rect 2791 24454 2805 24506
rect 2829 24454 2843 24506
rect 2843 24454 2855 24506
rect 2855 24454 2885 24506
rect 2909 24454 2919 24506
rect 2919 24454 2965 24506
rect 2669 24452 2725 24454
rect 2749 24452 2805 24454
rect 2829 24452 2885 24454
rect 2909 24452 2965 24454
rect 6096 24506 6152 24508
rect 6176 24506 6232 24508
rect 6256 24506 6312 24508
rect 6336 24506 6392 24508
rect 6096 24454 6142 24506
rect 6142 24454 6152 24506
rect 6176 24454 6206 24506
rect 6206 24454 6218 24506
rect 6218 24454 6232 24506
rect 6256 24454 6270 24506
rect 6270 24454 6282 24506
rect 6282 24454 6312 24506
rect 6336 24454 6346 24506
rect 6346 24454 6392 24506
rect 6096 24452 6152 24454
rect 6176 24452 6232 24454
rect 6256 24452 6312 24454
rect 6336 24452 6392 24454
rect 9523 24506 9579 24508
rect 9603 24506 9659 24508
rect 9683 24506 9739 24508
rect 9763 24506 9819 24508
rect 9523 24454 9569 24506
rect 9569 24454 9579 24506
rect 9603 24454 9633 24506
rect 9633 24454 9645 24506
rect 9645 24454 9659 24506
rect 9683 24454 9697 24506
rect 9697 24454 9709 24506
rect 9709 24454 9739 24506
rect 9763 24454 9773 24506
rect 9773 24454 9819 24506
rect 9523 24452 9579 24454
rect 9603 24452 9659 24454
rect 9683 24452 9739 24454
rect 9763 24452 9819 24454
rect 12950 24506 13006 24508
rect 13030 24506 13086 24508
rect 13110 24506 13166 24508
rect 13190 24506 13246 24508
rect 12950 24454 12996 24506
rect 12996 24454 13006 24506
rect 13030 24454 13060 24506
rect 13060 24454 13072 24506
rect 13072 24454 13086 24506
rect 13110 24454 13124 24506
rect 13124 24454 13136 24506
rect 13136 24454 13166 24506
rect 13190 24454 13200 24506
rect 13200 24454 13246 24506
rect 12950 24452 13006 24454
rect 13030 24452 13086 24454
rect 13110 24452 13166 24454
rect 13190 24452 13246 24454
rect 4382 23962 4438 23964
rect 4462 23962 4518 23964
rect 4542 23962 4598 23964
rect 4622 23962 4678 23964
rect 4382 23910 4428 23962
rect 4428 23910 4438 23962
rect 4462 23910 4492 23962
rect 4492 23910 4504 23962
rect 4504 23910 4518 23962
rect 4542 23910 4556 23962
rect 4556 23910 4568 23962
rect 4568 23910 4598 23962
rect 4622 23910 4632 23962
rect 4632 23910 4678 23962
rect 4382 23908 4438 23910
rect 4462 23908 4518 23910
rect 4542 23908 4598 23910
rect 4622 23908 4678 23910
rect 7809 23962 7865 23964
rect 7889 23962 7945 23964
rect 7969 23962 8025 23964
rect 8049 23962 8105 23964
rect 7809 23910 7855 23962
rect 7855 23910 7865 23962
rect 7889 23910 7919 23962
rect 7919 23910 7931 23962
rect 7931 23910 7945 23962
rect 7969 23910 7983 23962
rect 7983 23910 7995 23962
rect 7995 23910 8025 23962
rect 8049 23910 8059 23962
rect 8059 23910 8105 23962
rect 7809 23908 7865 23910
rect 7889 23908 7945 23910
rect 7969 23908 8025 23910
rect 8049 23908 8105 23910
rect 11236 23962 11292 23964
rect 11316 23962 11372 23964
rect 11396 23962 11452 23964
rect 11476 23962 11532 23964
rect 11236 23910 11282 23962
rect 11282 23910 11292 23962
rect 11316 23910 11346 23962
rect 11346 23910 11358 23962
rect 11358 23910 11372 23962
rect 11396 23910 11410 23962
rect 11410 23910 11422 23962
rect 11422 23910 11452 23962
rect 11476 23910 11486 23962
rect 11486 23910 11532 23962
rect 11236 23908 11292 23910
rect 11316 23908 11372 23910
rect 11396 23908 11452 23910
rect 11476 23908 11532 23910
rect 14663 23962 14719 23964
rect 14743 23962 14799 23964
rect 14823 23962 14879 23964
rect 14903 23962 14959 23964
rect 14663 23910 14709 23962
rect 14709 23910 14719 23962
rect 14743 23910 14773 23962
rect 14773 23910 14785 23962
rect 14785 23910 14799 23962
rect 14823 23910 14837 23962
rect 14837 23910 14849 23962
rect 14849 23910 14879 23962
rect 14903 23910 14913 23962
rect 14913 23910 14959 23962
rect 14663 23908 14719 23910
rect 14743 23908 14799 23910
rect 14823 23908 14879 23910
rect 14903 23908 14959 23910
rect 2669 23418 2725 23420
rect 2749 23418 2805 23420
rect 2829 23418 2885 23420
rect 2909 23418 2965 23420
rect 2669 23366 2715 23418
rect 2715 23366 2725 23418
rect 2749 23366 2779 23418
rect 2779 23366 2791 23418
rect 2791 23366 2805 23418
rect 2829 23366 2843 23418
rect 2843 23366 2855 23418
rect 2855 23366 2885 23418
rect 2909 23366 2919 23418
rect 2919 23366 2965 23418
rect 2669 23364 2725 23366
rect 2749 23364 2805 23366
rect 2829 23364 2885 23366
rect 2909 23364 2965 23366
rect 6096 23418 6152 23420
rect 6176 23418 6232 23420
rect 6256 23418 6312 23420
rect 6336 23418 6392 23420
rect 6096 23366 6142 23418
rect 6142 23366 6152 23418
rect 6176 23366 6206 23418
rect 6206 23366 6218 23418
rect 6218 23366 6232 23418
rect 6256 23366 6270 23418
rect 6270 23366 6282 23418
rect 6282 23366 6312 23418
rect 6336 23366 6346 23418
rect 6346 23366 6392 23418
rect 6096 23364 6152 23366
rect 6176 23364 6232 23366
rect 6256 23364 6312 23366
rect 6336 23364 6392 23366
rect 9523 23418 9579 23420
rect 9603 23418 9659 23420
rect 9683 23418 9739 23420
rect 9763 23418 9819 23420
rect 9523 23366 9569 23418
rect 9569 23366 9579 23418
rect 9603 23366 9633 23418
rect 9633 23366 9645 23418
rect 9645 23366 9659 23418
rect 9683 23366 9697 23418
rect 9697 23366 9709 23418
rect 9709 23366 9739 23418
rect 9763 23366 9773 23418
rect 9773 23366 9819 23418
rect 9523 23364 9579 23366
rect 9603 23364 9659 23366
rect 9683 23364 9739 23366
rect 9763 23364 9819 23366
rect 12950 23418 13006 23420
rect 13030 23418 13086 23420
rect 13110 23418 13166 23420
rect 13190 23418 13246 23420
rect 12950 23366 12996 23418
rect 12996 23366 13006 23418
rect 13030 23366 13060 23418
rect 13060 23366 13072 23418
rect 13072 23366 13086 23418
rect 13110 23366 13124 23418
rect 13124 23366 13136 23418
rect 13136 23366 13166 23418
rect 13190 23366 13200 23418
rect 13200 23366 13246 23418
rect 12950 23364 13006 23366
rect 13030 23364 13086 23366
rect 13110 23364 13166 23366
rect 13190 23364 13246 23366
rect 4382 22874 4438 22876
rect 4462 22874 4518 22876
rect 4542 22874 4598 22876
rect 4622 22874 4678 22876
rect 4382 22822 4428 22874
rect 4428 22822 4438 22874
rect 4462 22822 4492 22874
rect 4492 22822 4504 22874
rect 4504 22822 4518 22874
rect 4542 22822 4556 22874
rect 4556 22822 4568 22874
rect 4568 22822 4598 22874
rect 4622 22822 4632 22874
rect 4632 22822 4678 22874
rect 4382 22820 4438 22822
rect 4462 22820 4518 22822
rect 4542 22820 4598 22822
rect 4622 22820 4678 22822
rect 7809 22874 7865 22876
rect 7889 22874 7945 22876
rect 7969 22874 8025 22876
rect 8049 22874 8105 22876
rect 7809 22822 7855 22874
rect 7855 22822 7865 22874
rect 7889 22822 7919 22874
rect 7919 22822 7931 22874
rect 7931 22822 7945 22874
rect 7969 22822 7983 22874
rect 7983 22822 7995 22874
rect 7995 22822 8025 22874
rect 8049 22822 8059 22874
rect 8059 22822 8105 22874
rect 7809 22820 7865 22822
rect 7889 22820 7945 22822
rect 7969 22820 8025 22822
rect 8049 22820 8105 22822
rect 11236 22874 11292 22876
rect 11316 22874 11372 22876
rect 11396 22874 11452 22876
rect 11476 22874 11532 22876
rect 11236 22822 11282 22874
rect 11282 22822 11292 22874
rect 11316 22822 11346 22874
rect 11346 22822 11358 22874
rect 11358 22822 11372 22874
rect 11396 22822 11410 22874
rect 11410 22822 11422 22874
rect 11422 22822 11452 22874
rect 11476 22822 11486 22874
rect 11486 22822 11532 22874
rect 11236 22820 11292 22822
rect 11316 22820 11372 22822
rect 11396 22820 11452 22822
rect 11476 22820 11532 22822
rect 14663 22874 14719 22876
rect 14743 22874 14799 22876
rect 14823 22874 14879 22876
rect 14903 22874 14959 22876
rect 14663 22822 14709 22874
rect 14709 22822 14719 22874
rect 14743 22822 14773 22874
rect 14773 22822 14785 22874
rect 14785 22822 14799 22874
rect 14823 22822 14837 22874
rect 14837 22822 14849 22874
rect 14849 22822 14879 22874
rect 14903 22822 14913 22874
rect 14913 22822 14959 22874
rect 14663 22820 14719 22822
rect 14743 22820 14799 22822
rect 14823 22820 14879 22822
rect 14903 22820 14959 22822
rect 2669 22330 2725 22332
rect 2749 22330 2805 22332
rect 2829 22330 2885 22332
rect 2909 22330 2965 22332
rect 2669 22278 2715 22330
rect 2715 22278 2725 22330
rect 2749 22278 2779 22330
rect 2779 22278 2791 22330
rect 2791 22278 2805 22330
rect 2829 22278 2843 22330
rect 2843 22278 2855 22330
rect 2855 22278 2885 22330
rect 2909 22278 2919 22330
rect 2919 22278 2965 22330
rect 2669 22276 2725 22278
rect 2749 22276 2805 22278
rect 2829 22276 2885 22278
rect 2909 22276 2965 22278
rect 6096 22330 6152 22332
rect 6176 22330 6232 22332
rect 6256 22330 6312 22332
rect 6336 22330 6392 22332
rect 6096 22278 6142 22330
rect 6142 22278 6152 22330
rect 6176 22278 6206 22330
rect 6206 22278 6218 22330
rect 6218 22278 6232 22330
rect 6256 22278 6270 22330
rect 6270 22278 6282 22330
rect 6282 22278 6312 22330
rect 6336 22278 6346 22330
rect 6346 22278 6392 22330
rect 6096 22276 6152 22278
rect 6176 22276 6232 22278
rect 6256 22276 6312 22278
rect 6336 22276 6392 22278
rect 9523 22330 9579 22332
rect 9603 22330 9659 22332
rect 9683 22330 9739 22332
rect 9763 22330 9819 22332
rect 9523 22278 9569 22330
rect 9569 22278 9579 22330
rect 9603 22278 9633 22330
rect 9633 22278 9645 22330
rect 9645 22278 9659 22330
rect 9683 22278 9697 22330
rect 9697 22278 9709 22330
rect 9709 22278 9739 22330
rect 9763 22278 9773 22330
rect 9773 22278 9819 22330
rect 9523 22276 9579 22278
rect 9603 22276 9659 22278
rect 9683 22276 9739 22278
rect 9763 22276 9819 22278
rect 12950 22330 13006 22332
rect 13030 22330 13086 22332
rect 13110 22330 13166 22332
rect 13190 22330 13246 22332
rect 12950 22278 12996 22330
rect 12996 22278 13006 22330
rect 13030 22278 13060 22330
rect 13060 22278 13072 22330
rect 13072 22278 13086 22330
rect 13110 22278 13124 22330
rect 13124 22278 13136 22330
rect 13136 22278 13166 22330
rect 13190 22278 13200 22330
rect 13200 22278 13246 22330
rect 12950 22276 13006 22278
rect 13030 22276 13086 22278
rect 13110 22276 13166 22278
rect 13190 22276 13246 22278
rect 4382 21786 4438 21788
rect 4462 21786 4518 21788
rect 4542 21786 4598 21788
rect 4622 21786 4678 21788
rect 4382 21734 4428 21786
rect 4428 21734 4438 21786
rect 4462 21734 4492 21786
rect 4492 21734 4504 21786
rect 4504 21734 4518 21786
rect 4542 21734 4556 21786
rect 4556 21734 4568 21786
rect 4568 21734 4598 21786
rect 4622 21734 4632 21786
rect 4632 21734 4678 21786
rect 4382 21732 4438 21734
rect 4462 21732 4518 21734
rect 4542 21732 4598 21734
rect 4622 21732 4678 21734
rect 7809 21786 7865 21788
rect 7889 21786 7945 21788
rect 7969 21786 8025 21788
rect 8049 21786 8105 21788
rect 7809 21734 7855 21786
rect 7855 21734 7865 21786
rect 7889 21734 7919 21786
rect 7919 21734 7931 21786
rect 7931 21734 7945 21786
rect 7969 21734 7983 21786
rect 7983 21734 7995 21786
rect 7995 21734 8025 21786
rect 8049 21734 8059 21786
rect 8059 21734 8105 21786
rect 7809 21732 7865 21734
rect 7889 21732 7945 21734
rect 7969 21732 8025 21734
rect 8049 21732 8105 21734
rect 11236 21786 11292 21788
rect 11316 21786 11372 21788
rect 11396 21786 11452 21788
rect 11476 21786 11532 21788
rect 11236 21734 11282 21786
rect 11282 21734 11292 21786
rect 11316 21734 11346 21786
rect 11346 21734 11358 21786
rect 11358 21734 11372 21786
rect 11396 21734 11410 21786
rect 11410 21734 11422 21786
rect 11422 21734 11452 21786
rect 11476 21734 11486 21786
rect 11486 21734 11532 21786
rect 11236 21732 11292 21734
rect 11316 21732 11372 21734
rect 11396 21732 11452 21734
rect 11476 21732 11532 21734
rect 14663 21786 14719 21788
rect 14743 21786 14799 21788
rect 14823 21786 14879 21788
rect 14903 21786 14959 21788
rect 14663 21734 14709 21786
rect 14709 21734 14719 21786
rect 14743 21734 14773 21786
rect 14773 21734 14785 21786
rect 14785 21734 14799 21786
rect 14823 21734 14837 21786
rect 14837 21734 14849 21786
rect 14849 21734 14879 21786
rect 14903 21734 14913 21786
rect 14913 21734 14959 21786
rect 14663 21732 14719 21734
rect 14743 21732 14799 21734
rect 14823 21732 14879 21734
rect 14903 21732 14959 21734
rect 2669 21242 2725 21244
rect 2749 21242 2805 21244
rect 2829 21242 2885 21244
rect 2909 21242 2965 21244
rect 2669 21190 2715 21242
rect 2715 21190 2725 21242
rect 2749 21190 2779 21242
rect 2779 21190 2791 21242
rect 2791 21190 2805 21242
rect 2829 21190 2843 21242
rect 2843 21190 2855 21242
rect 2855 21190 2885 21242
rect 2909 21190 2919 21242
rect 2919 21190 2965 21242
rect 2669 21188 2725 21190
rect 2749 21188 2805 21190
rect 2829 21188 2885 21190
rect 2909 21188 2965 21190
rect 6096 21242 6152 21244
rect 6176 21242 6232 21244
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6096 21190 6142 21242
rect 6142 21190 6152 21242
rect 6176 21190 6206 21242
rect 6206 21190 6218 21242
rect 6218 21190 6232 21242
rect 6256 21190 6270 21242
rect 6270 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6096 21188 6152 21190
rect 6176 21188 6232 21190
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 9523 21242 9579 21244
rect 9603 21242 9659 21244
rect 9683 21242 9739 21244
rect 9763 21242 9819 21244
rect 9523 21190 9569 21242
rect 9569 21190 9579 21242
rect 9603 21190 9633 21242
rect 9633 21190 9645 21242
rect 9645 21190 9659 21242
rect 9683 21190 9697 21242
rect 9697 21190 9709 21242
rect 9709 21190 9739 21242
rect 9763 21190 9773 21242
rect 9773 21190 9819 21242
rect 9523 21188 9579 21190
rect 9603 21188 9659 21190
rect 9683 21188 9739 21190
rect 9763 21188 9819 21190
rect 12950 21242 13006 21244
rect 13030 21242 13086 21244
rect 13110 21242 13166 21244
rect 13190 21242 13246 21244
rect 12950 21190 12996 21242
rect 12996 21190 13006 21242
rect 13030 21190 13060 21242
rect 13060 21190 13072 21242
rect 13072 21190 13086 21242
rect 13110 21190 13124 21242
rect 13124 21190 13136 21242
rect 13136 21190 13166 21242
rect 13190 21190 13200 21242
rect 13200 21190 13246 21242
rect 12950 21188 13006 21190
rect 13030 21188 13086 21190
rect 13110 21188 13166 21190
rect 13190 21188 13246 21190
rect 4382 20698 4438 20700
rect 4462 20698 4518 20700
rect 4542 20698 4598 20700
rect 4622 20698 4678 20700
rect 4382 20646 4428 20698
rect 4428 20646 4438 20698
rect 4462 20646 4492 20698
rect 4492 20646 4504 20698
rect 4504 20646 4518 20698
rect 4542 20646 4556 20698
rect 4556 20646 4568 20698
rect 4568 20646 4598 20698
rect 4622 20646 4632 20698
rect 4632 20646 4678 20698
rect 4382 20644 4438 20646
rect 4462 20644 4518 20646
rect 4542 20644 4598 20646
rect 4622 20644 4678 20646
rect 7809 20698 7865 20700
rect 7889 20698 7945 20700
rect 7969 20698 8025 20700
rect 8049 20698 8105 20700
rect 7809 20646 7855 20698
rect 7855 20646 7865 20698
rect 7889 20646 7919 20698
rect 7919 20646 7931 20698
rect 7931 20646 7945 20698
rect 7969 20646 7983 20698
rect 7983 20646 7995 20698
rect 7995 20646 8025 20698
rect 8049 20646 8059 20698
rect 8059 20646 8105 20698
rect 7809 20644 7865 20646
rect 7889 20644 7945 20646
rect 7969 20644 8025 20646
rect 8049 20644 8105 20646
rect 11236 20698 11292 20700
rect 11316 20698 11372 20700
rect 11396 20698 11452 20700
rect 11476 20698 11532 20700
rect 11236 20646 11282 20698
rect 11282 20646 11292 20698
rect 11316 20646 11346 20698
rect 11346 20646 11358 20698
rect 11358 20646 11372 20698
rect 11396 20646 11410 20698
rect 11410 20646 11422 20698
rect 11422 20646 11452 20698
rect 11476 20646 11486 20698
rect 11486 20646 11532 20698
rect 11236 20644 11292 20646
rect 11316 20644 11372 20646
rect 11396 20644 11452 20646
rect 11476 20644 11532 20646
rect 14663 20698 14719 20700
rect 14743 20698 14799 20700
rect 14823 20698 14879 20700
rect 14903 20698 14959 20700
rect 14663 20646 14709 20698
rect 14709 20646 14719 20698
rect 14743 20646 14773 20698
rect 14773 20646 14785 20698
rect 14785 20646 14799 20698
rect 14823 20646 14837 20698
rect 14837 20646 14849 20698
rect 14849 20646 14879 20698
rect 14903 20646 14913 20698
rect 14913 20646 14959 20698
rect 14663 20644 14719 20646
rect 14743 20644 14799 20646
rect 14823 20644 14879 20646
rect 14903 20644 14959 20646
rect 2669 20154 2725 20156
rect 2749 20154 2805 20156
rect 2829 20154 2885 20156
rect 2909 20154 2965 20156
rect 2669 20102 2715 20154
rect 2715 20102 2725 20154
rect 2749 20102 2779 20154
rect 2779 20102 2791 20154
rect 2791 20102 2805 20154
rect 2829 20102 2843 20154
rect 2843 20102 2855 20154
rect 2855 20102 2885 20154
rect 2909 20102 2919 20154
rect 2919 20102 2965 20154
rect 2669 20100 2725 20102
rect 2749 20100 2805 20102
rect 2829 20100 2885 20102
rect 2909 20100 2965 20102
rect 6096 20154 6152 20156
rect 6176 20154 6232 20156
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6096 20102 6142 20154
rect 6142 20102 6152 20154
rect 6176 20102 6206 20154
rect 6206 20102 6218 20154
rect 6218 20102 6232 20154
rect 6256 20102 6270 20154
rect 6270 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6096 20100 6152 20102
rect 6176 20100 6232 20102
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 9523 20154 9579 20156
rect 9603 20154 9659 20156
rect 9683 20154 9739 20156
rect 9763 20154 9819 20156
rect 9523 20102 9569 20154
rect 9569 20102 9579 20154
rect 9603 20102 9633 20154
rect 9633 20102 9645 20154
rect 9645 20102 9659 20154
rect 9683 20102 9697 20154
rect 9697 20102 9709 20154
rect 9709 20102 9739 20154
rect 9763 20102 9773 20154
rect 9773 20102 9819 20154
rect 9523 20100 9579 20102
rect 9603 20100 9659 20102
rect 9683 20100 9739 20102
rect 9763 20100 9819 20102
rect 12950 20154 13006 20156
rect 13030 20154 13086 20156
rect 13110 20154 13166 20156
rect 13190 20154 13246 20156
rect 12950 20102 12996 20154
rect 12996 20102 13006 20154
rect 13030 20102 13060 20154
rect 13060 20102 13072 20154
rect 13072 20102 13086 20154
rect 13110 20102 13124 20154
rect 13124 20102 13136 20154
rect 13136 20102 13166 20154
rect 13190 20102 13200 20154
rect 13200 20102 13246 20154
rect 12950 20100 13006 20102
rect 13030 20100 13086 20102
rect 13110 20100 13166 20102
rect 13190 20100 13246 20102
rect 14462 19896 14518 19952
rect 4382 19610 4438 19612
rect 4462 19610 4518 19612
rect 4542 19610 4598 19612
rect 4622 19610 4678 19612
rect 4382 19558 4428 19610
rect 4428 19558 4438 19610
rect 4462 19558 4492 19610
rect 4492 19558 4504 19610
rect 4504 19558 4518 19610
rect 4542 19558 4556 19610
rect 4556 19558 4568 19610
rect 4568 19558 4598 19610
rect 4622 19558 4632 19610
rect 4632 19558 4678 19610
rect 4382 19556 4438 19558
rect 4462 19556 4518 19558
rect 4542 19556 4598 19558
rect 4622 19556 4678 19558
rect 7809 19610 7865 19612
rect 7889 19610 7945 19612
rect 7969 19610 8025 19612
rect 8049 19610 8105 19612
rect 7809 19558 7855 19610
rect 7855 19558 7865 19610
rect 7889 19558 7919 19610
rect 7919 19558 7931 19610
rect 7931 19558 7945 19610
rect 7969 19558 7983 19610
rect 7983 19558 7995 19610
rect 7995 19558 8025 19610
rect 8049 19558 8059 19610
rect 8059 19558 8105 19610
rect 7809 19556 7865 19558
rect 7889 19556 7945 19558
rect 7969 19556 8025 19558
rect 8049 19556 8105 19558
rect 11236 19610 11292 19612
rect 11316 19610 11372 19612
rect 11396 19610 11452 19612
rect 11476 19610 11532 19612
rect 11236 19558 11282 19610
rect 11282 19558 11292 19610
rect 11316 19558 11346 19610
rect 11346 19558 11358 19610
rect 11358 19558 11372 19610
rect 11396 19558 11410 19610
rect 11410 19558 11422 19610
rect 11422 19558 11452 19610
rect 11476 19558 11486 19610
rect 11486 19558 11532 19610
rect 11236 19556 11292 19558
rect 11316 19556 11372 19558
rect 11396 19556 11452 19558
rect 11476 19556 11532 19558
rect 14663 19610 14719 19612
rect 14743 19610 14799 19612
rect 14823 19610 14879 19612
rect 14903 19610 14959 19612
rect 14663 19558 14709 19610
rect 14709 19558 14719 19610
rect 14743 19558 14773 19610
rect 14773 19558 14785 19610
rect 14785 19558 14799 19610
rect 14823 19558 14837 19610
rect 14837 19558 14849 19610
rect 14849 19558 14879 19610
rect 14903 19558 14913 19610
rect 14913 19558 14959 19610
rect 14663 19556 14719 19558
rect 14743 19556 14799 19558
rect 14823 19556 14879 19558
rect 14903 19556 14959 19558
rect 2669 19066 2725 19068
rect 2749 19066 2805 19068
rect 2829 19066 2885 19068
rect 2909 19066 2965 19068
rect 2669 19014 2715 19066
rect 2715 19014 2725 19066
rect 2749 19014 2779 19066
rect 2779 19014 2791 19066
rect 2791 19014 2805 19066
rect 2829 19014 2843 19066
rect 2843 19014 2855 19066
rect 2855 19014 2885 19066
rect 2909 19014 2919 19066
rect 2919 19014 2965 19066
rect 2669 19012 2725 19014
rect 2749 19012 2805 19014
rect 2829 19012 2885 19014
rect 2909 19012 2965 19014
rect 6096 19066 6152 19068
rect 6176 19066 6232 19068
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6096 19014 6142 19066
rect 6142 19014 6152 19066
rect 6176 19014 6206 19066
rect 6206 19014 6218 19066
rect 6218 19014 6232 19066
rect 6256 19014 6270 19066
rect 6270 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6096 19012 6152 19014
rect 6176 19012 6232 19014
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 9523 19066 9579 19068
rect 9603 19066 9659 19068
rect 9683 19066 9739 19068
rect 9763 19066 9819 19068
rect 9523 19014 9569 19066
rect 9569 19014 9579 19066
rect 9603 19014 9633 19066
rect 9633 19014 9645 19066
rect 9645 19014 9659 19066
rect 9683 19014 9697 19066
rect 9697 19014 9709 19066
rect 9709 19014 9739 19066
rect 9763 19014 9773 19066
rect 9773 19014 9819 19066
rect 9523 19012 9579 19014
rect 9603 19012 9659 19014
rect 9683 19012 9739 19014
rect 9763 19012 9819 19014
rect 12950 19066 13006 19068
rect 13030 19066 13086 19068
rect 13110 19066 13166 19068
rect 13190 19066 13246 19068
rect 12950 19014 12996 19066
rect 12996 19014 13006 19066
rect 13030 19014 13060 19066
rect 13060 19014 13072 19066
rect 13072 19014 13086 19066
rect 13110 19014 13124 19066
rect 13124 19014 13136 19066
rect 13136 19014 13166 19066
rect 13190 19014 13200 19066
rect 13200 19014 13246 19066
rect 12950 19012 13006 19014
rect 13030 19012 13086 19014
rect 13110 19012 13166 19014
rect 13190 19012 13246 19014
rect 4382 18522 4438 18524
rect 4462 18522 4518 18524
rect 4542 18522 4598 18524
rect 4622 18522 4678 18524
rect 4382 18470 4428 18522
rect 4428 18470 4438 18522
rect 4462 18470 4492 18522
rect 4492 18470 4504 18522
rect 4504 18470 4518 18522
rect 4542 18470 4556 18522
rect 4556 18470 4568 18522
rect 4568 18470 4598 18522
rect 4622 18470 4632 18522
rect 4632 18470 4678 18522
rect 4382 18468 4438 18470
rect 4462 18468 4518 18470
rect 4542 18468 4598 18470
rect 4622 18468 4678 18470
rect 7809 18522 7865 18524
rect 7889 18522 7945 18524
rect 7969 18522 8025 18524
rect 8049 18522 8105 18524
rect 7809 18470 7855 18522
rect 7855 18470 7865 18522
rect 7889 18470 7919 18522
rect 7919 18470 7931 18522
rect 7931 18470 7945 18522
rect 7969 18470 7983 18522
rect 7983 18470 7995 18522
rect 7995 18470 8025 18522
rect 8049 18470 8059 18522
rect 8059 18470 8105 18522
rect 7809 18468 7865 18470
rect 7889 18468 7945 18470
rect 7969 18468 8025 18470
rect 8049 18468 8105 18470
rect 11236 18522 11292 18524
rect 11316 18522 11372 18524
rect 11396 18522 11452 18524
rect 11476 18522 11532 18524
rect 11236 18470 11282 18522
rect 11282 18470 11292 18522
rect 11316 18470 11346 18522
rect 11346 18470 11358 18522
rect 11358 18470 11372 18522
rect 11396 18470 11410 18522
rect 11410 18470 11422 18522
rect 11422 18470 11452 18522
rect 11476 18470 11486 18522
rect 11486 18470 11532 18522
rect 11236 18468 11292 18470
rect 11316 18468 11372 18470
rect 11396 18468 11452 18470
rect 11476 18468 11532 18470
rect 14663 18522 14719 18524
rect 14743 18522 14799 18524
rect 14823 18522 14879 18524
rect 14903 18522 14959 18524
rect 14663 18470 14709 18522
rect 14709 18470 14719 18522
rect 14743 18470 14773 18522
rect 14773 18470 14785 18522
rect 14785 18470 14799 18522
rect 14823 18470 14837 18522
rect 14837 18470 14849 18522
rect 14849 18470 14879 18522
rect 14903 18470 14913 18522
rect 14913 18470 14959 18522
rect 14663 18468 14719 18470
rect 14743 18468 14799 18470
rect 14823 18468 14879 18470
rect 14903 18468 14959 18470
rect 2669 17978 2725 17980
rect 2749 17978 2805 17980
rect 2829 17978 2885 17980
rect 2909 17978 2965 17980
rect 2669 17926 2715 17978
rect 2715 17926 2725 17978
rect 2749 17926 2779 17978
rect 2779 17926 2791 17978
rect 2791 17926 2805 17978
rect 2829 17926 2843 17978
rect 2843 17926 2855 17978
rect 2855 17926 2885 17978
rect 2909 17926 2919 17978
rect 2919 17926 2965 17978
rect 2669 17924 2725 17926
rect 2749 17924 2805 17926
rect 2829 17924 2885 17926
rect 2909 17924 2965 17926
rect 6096 17978 6152 17980
rect 6176 17978 6232 17980
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6096 17926 6142 17978
rect 6142 17926 6152 17978
rect 6176 17926 6206 17978
rect 6206 17926 6218 17978
rect 6218 17926 6232 17978
rect 6256 17926 6270 17978
rect 6270 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6096 17924 6152 17926
rect 6176 17924 6232 17926
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 9523 17978 9579 17980
rect 9603 17978 9659 17980
rect 9683 17978 9739 17980
rect 9763 17978 9819 17980
rect 9523 17926 9569 17978
rect 9569 17926 9579 17978
rect 9603 17926 9633 17978
rect 9633 17926 9645 17978
rect 9645 17926 9659 17978
rect 9683 17926 9697 17978
rect 9697 17926 9709 17978
rect 9709 17926 9739 17978
rect 9763 17926 9773 17978
rect 9773 17926 9819 17978
rect 9523 17924 9579 17926
rect 9603 17924 9659 17926
rect 9683 17924 9739 17926
rect 9763 17924 9819 17926
rect 12950 17978 13006 17980
rect 13030 17978 13086 17980
rect 13110 17978 13166 17980
rect 13190 17978 13246 17980
rect 12950 17926 12996 17978
rect 12996 17926 13006 17978
rect 13030 17926 13060 17978
rect 13060 17926 13072 17978
rect 13072 17926 13086 17978
rect 13110 17926 13124 17978
rect 13124 17926 13136 17978
rect 13136 17926 13166 17978
rect 13190 17926 13200 17978
rect 13200 17926 13246 17978
rect 12950 17924 13006 17926
rect 13030 17924 13086 17926
rect 13110 17924 13166 17926
rect 13190 17924 13246 17926
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 14462 12164 14518 12200
rect 14462 12144 14464 12164
rect 14464 12144 14516 12164
rect 14516 12144 14518 12164
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14462 4120 14518 4176
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
<< metal3 >>
rect 4372 45728 4688 45729
rect 4372 45664 4378 45728
rect 4442 45664 4458 45728
rect 4522 45664 4538 45728
rect 4602 45664 4618 45728
rect 4682 45664 4688 45728
rect 4372 45663 4688 45664
rect 7799 45728 8115 45729
rect 7799 45664 7805 45728
rect 7869 45664 7885 45728
rect 7949 45664 7965 45728
rect 8029 45664 8045 45728
rect 8109 45664 8115 45728
rect 7799 45663 8115 45664
rect 11226 45728 11542 45729
rect 11226 45664 11232 45728
rect 11296 45664 11312 45728
rect 11376 45664 11392 45728
rect 11456 45664 11472 45728
rect 11536 45664 11542 45728
rect 11226 45663 11542 45664
rect 14653 45728 14969 45729
rect 14653 45664 14659 45728
rect 14723 45664 14739 45728
rect 14803 45664 14819 45728
rect 14883 45664 14899 45728
rect 14963 45664 14969 45728
rect 14653 45663 14969 45664
rect 2659 45184 2975 45185
rect 2659 45120 2665 45184
rect 2729 45120 2745 45184
rect 2809 45120 2825 45184
rect 2889 45120 2905 45184
rect 2969 45120 2975 45184
rect 2659 45119 2975 45120
rect 6086 45184 6402 45185
rect 6086 45120 6092 45184
rect 6156 45120 6172 45184
rect 6236 45120 6252 45184
rect 6316 45120 6332 45184
rect 6396 45120 6402 45184
rect 6086 45119 6402 45120
rect 9513 45184 9829 45185
rect 9513 45120 9519 45184
rect 9583 45120 9599 45184
rect 9663 45120 9679 45184
rect 9743 45120 9759 45184
rect 9823 45120 9829 45184
rect 9513 45119 9829 45120
rect 12940 45184 13256 45185
rect 12940 45120 12946 45184
rect 13010 45120 13026 45184
rect 13090 45120 13106 45184
rect 13170 45120 13186 45184
rect 13250 45120 13256 45184
rect 12940 45119 13256 45120
rect 4372 44640 4688 44641
rect 4372 44576 4378 44640
rect 4442 44576 4458 44640
rect 4522 44576 4538 44640
rect 4602 44576 4618 44640
rect 4682 44576 4688 44640
rect 4372 44575 4688 44576
rect 7799 44640 8115 44641
rect 7799 44576 7805 44640
rect 7869 44576 7885 44640
rect 7949 44576 7965 44640
rect 8029 44576 8045 44640
rect 8109 44576 8115 44640
rect 7799 44575 8115 44576
rect 11226 44640 11542 44641
rect 11226 44576 11232 44640
rect 11296 44576 11312 44640
rect 11376 44576 11392 44640
rect 11456 44576 11472 44640
rect 11536 44576 11542 44640
rect 11226 44575 11542 44576
rect 14653 44640 14969 44641
rect 14653 44576 14659 44640
rect 14723 44576 14739 44640
rect 14803 44576 14819 44640
rect 14883 44576 14899 44640
rect 14963 44576 14969 44640
rect 14653 44575 14969 44576
rect 2659 44096 2975 44097
rect 2659 44032 2665 44096
rect 2729 44032 2745 44096
rect 2809 44032 2825 44096
rect 2889 44032 2905 44096
rect 2969 44032 2975 44096
rect 2659 44031 2975 44032
rect 6086 44096 6402 44097
rect 6086 44032 6092 44096
rect 6156 44032 6172 44096
rect 6236 44032 6252 44096
rect 6316 44032 6332 44096
rect 6396 44032 6402 44096
rect 6086 44031 6402 44032
rect 9513 44096 9829 44097
rect 9513 44032 9519 44096
rect 9583 44032 9599 44096
rect 9663 44032 9679 44096
rect 9743 44032 9759 44096
rect 9823 44032 9829 44096
rect 9513 44031 9829 44032
rect 12940 44096 13256 44097
rect 12940 44032 12946 44096
rect 13010 44032 13026 44096
rect 13090 44032 13106 44096
rect 13170 44032 13186 44096
rect 13250 44032 13256 44096
rect 12940 44031 13256 44032
rect 14457 43754 14523 43757
rect 14457 43752 15210 43754
rect 14457 43696 14462 43752
rect 14518 43696 15210 43752
rect 14457 43694 15210 43696
rect 14457 43691 14523 43694
rect 15150 43648 15210 43694
rect 15150 43558 16000 43648
rect 4372 43552 4688 43553
rect 4372 43488 4378 43552
rect 4442 43488 4458 43552
rect 4522 43488 4538 43552
rect 4602 43488 4618 43552
rect 4682 43488 4688 43552
rect 4372 43487 4688 43488
rect 7799 43552 8115 43553
rect 7799 43488 7805 43552
rect 7869 43488 7885 43552
rect 7949 43488 7965 43552
rect 8029 43488 8045 43552
rect 8109 43488 8115 43552
rect 7799 43487 8115 43488
rect 11226 43552 11542 43553
rect 11226 43488 11232 43552
rect 11296 43488 11312 43552
rect 11376 43488 11392 43552
rect 11456 43488 11472 43552
rect 11536 43488 11542 43552
rect 11226 43487 11542 43488
rect 14653 43552 14969 43553
rect 14653 43488 14659 43552
rect 14723 43488 14739 43552
rect 14803 43488 14819 43552
rect 14883 43488 14899 43552
rect 14963 43488 14969 43552
rect 15200 43528 16000 43558
rect 14653 43487 14969 43488
rect 2659 43008 2975 43009
rect 2659 42944 2665 43008
rect 2729 42944 2745 43008
rect 2809 42944 2825 43008
rect 2889 42944 2905 43008
rect 2969 42944 2975 43008
rect 2659 42943 2975 42944
rect 6086 43008 6402 43009
rect 6086 42944 6092 43008
rect 6156 42944 6172 43008
rect 6236 42944 6252 43008
rect 6316 42944 6332 43008
rect 6396 42944 6402 43008
rect 6086 42943 6402 42944
rect 9513 43008 9829 43009
rect 9513 42944 9519 43008
rect 9583 42944 9599 43008
rect 9663 42944 9679 43008
rect 9743 42944 9759 43008
rect 9823 42944 9829 43008
rect 9513 42943 9829 42944
rect 12940 43008 13256 43009
rect 12940 42944 12946 43008
rect 13010 42944 13026 43008
rect 13090 42944 13106 43008
rect 13170 42944 13186 43008
rect 13250 42944 13256 43008
rect 12940 42943 13256 42944
rect 4372 42464 4688 42465
rect 4372 42400 4378 42464
rect 4442 42400 4458 42464
rect 4522 42400 4538 42464
rect 4602 42400 4618 42464
rect 4682 42400 4688 42464
rect 4372 42399 4688 42400
rect 7799 42464 8115 42465
rect 7799 42400 7805 42464
rect 7869 42400 7885 42464
rect 7949 42400 7965 42464
rect 8029 42400 8045 42464
rect 8109 42400 8115 42464
rect 7799 42399 8115 42400
rect 11226 42464 11542 42465
rect 11226 42400 11232 42464
rect 11296 42400 11312 42464
rect 11376 42400 11392 42464
rect 11456 42400 11472 42464
rect 11536 42400 11542 42464
rect 11226 42399 11542 42400
rect 14653 42464 14969 42465
rect 14653 42400 14659 42464
rect 14723 42400 14739 42464
rect 14803 42400 14819 42464
rect 14883 42400 14899 42464
rect 14963 42400 14969 42464
rect 14653 42399 14969 42400
rect 2659 41920 2975 41921
rect 2659 41856 2665 41920
rect 2729 41856 2745 41920
rect 2809 41856 2825 41920
rect 2889 41856 2905 41920
rect 2969 41856 2975 41920
rect 2659 41855 2975 41856
rect 6086 41920 6402 41921
rect 6086 41856 6092 41920
rect 6156 41856 6172 41920
rect 6236 41856 6252 41920
rect 6316 41856 6332 41920
rect 6396 41856 6402 41920
rect 6086 41855 6402 41856
rect 9513 41920 9829 41921
rect 9513 41856 9519 41920
rect 9583 41856 9599 41920
rect 9663 41856 9679 41920
rect 9743 41856 9759 41920
rect 9823 41856 9829 41920
rect 9513 41855 9829 41856
rect 12940 41920 13256 41921
rect 12940 41856 12946 41920
rect 13010 41856 13026 41920
rect 13090 41856 13106 41920
rect 13170 41856 13186 41920
rect 13250 41856 13256 41920
rect 12940 41855 13256 41856
rect 4372 41376 4688 41377
rect 4372 41312 4378 41376
rect 4442 41312 4458 41376
rect 4522 41312 4538 41376
rect 4602 41312 4618 41376
rect 4682 41312 4688 41376
rect 4372 41311 4688 41312
rect 7799 41376 8115 41377
rect 7799 41312 7805 41376
rect 7869 41312 7885 41376
rect 7949 41312 7965 41376
rect 8029 41312 8045 41376
rect 8109 41312 8115 41376
rect 7799 41311 8115 41312
rect 11226 41376 11542 41377
rect 11226 41312 11232 41376
rect 11296 41312 11312 41376
rect 11376 41312 11392 41376
rect 11456 41312 11472 41376
rect 11536 41312 11542 41376
rect 11226 41311 11542 41312
rect 14653 41376 14969 41377
rect 14653 41312 14659 41376
rect 14723 41312 14739 41376
rect 14803 41312 14819 41376
rect 14883 41312 14899 41376
rect 14963 41312 14969 41376
rect 14653 41311 14969 41312
rect 2659 40832 2975 40833
rect 2659 40768 2665 40832
rect 2729 40768 2745 40832
rect 2809 40768 2825 40832
rect 2889 40768 2905 40832
rect 2969 40768 2975 40832
rect 2659 40767 2975 40768
rect 6086 40832 6402 40833
rect 6086 40768 6092 40832
rect 6156 40768 6172 40832
rect 6236 40768 6252 40832
rect 6316 40768 6332 40832
rect 6396 40768 6402 40832
rect 6086 40767 6402 40768
rect 9513 40832 9829 40833
rect 9513 40768 9519 40832
rect 9583 40768 9599 40832
rect 9663 40768 9679 40832
rect 9743 40768 9759 40832
rect 9823 40768 9829 40832
rect 9513 40767 9829 40768
rect 12940 40832 13256 40833
rect 12940 40768 12946 40832
rect 13010 40768 13026 40832
rect 13090 40768 13106 40832
rect 13170 40768 13186 40832
rect 13250 40768 13256 40832
rect 12940 40767 13256 40768
rect 4372 40288 4688 40289
rect 4372 40224 4378 40288
rect 4442 40224 4458 40288
rect 4522 40224 4538 40288
rect 4602 40224 4618 40288
rect 4682 40224 4688 40288
rect 4372 40223 4688 40224
rect 7799 40288 8115 40289
rect 7799 40224 7805 40288
rect 7869 40224 7885 40288
rect 7949 40224 7965 40288
rect 8029 40224 8045 40288
rect 8109 40224 8115 40288
rect 7799 40223 8115 40224
rect 11226 40288 11542 40289
rect 11226 40224 11232 40288
rect 11296 40224 11312 40288
rect 11376 40224 11392 40288
rect 11456 40224 11472 40288
rect 11536 40224 11542 40288
rect 11226 40223 11542 40224
rect 14653 40288 14969 40289
rect 14653 40224 14659 40288
rect 14723 40224 14739 40288
rect 14803 40224 14819 40288
rect 14883 40224 14899 40288
rect 14963 40224 14969 40288
rect 14653 40223 14969 40224
rect 2659 39744 2975 39745
rect 2659 39680 2665 39744
rect 2729 39680 2745 39744
rect 2809 39680 2825 39744
rect 2889 39680 2905 39744
rect 2969 39680 2975 39744
rect 2659 39679 2975 39680
rect 6086 39744 6402 39745
rect 6086 39680 6092 39744
rect 6156 39680 6172 39744
rect 6236 39680 6252 39744
rect 6316 39680 6332 39744
rect 6396 39680 6402 39744
rect 6086 39679 6402 39680
rect 9513 39744 9829 39745
rect 9513 39680 9519 39744
rect 9583 39680 9599 39744
rect 9663 39680 9679 39744
rect 9743 39680 9759 39744
rect 9823 39680 9829 39744
rect 9513 39679 9829 39680
rect 12940 39744 13256 39745
rect 12940 39680 12946 39744
rect 13010 39680 13026 39744
rect 13090 39680 13106 39744
rect 13170 39680 13186 39744
rect 13250 39680 13256 39744
rect 12940 39679 13256 39680
rect 4372 39200 4688 39201
rect 4372 39136 4378 39200
rect 4442 39136 4458 39200
rect 4522 39136 4538 39200
rect 4602 39136 4618 39200
rect 4682 39136 4688 39200
rect 4372 39135 4688 39136
rect 7799 39200 8115 39201
rect 7799 39136 7805 39200
rect 7869 39136 7885 39200
rect 7949 39136 7965 39200
rect 8029 39136 8045 39200
rect 8109 39136 8115 39200
rect 7799 39135 8115 39136
rect 11226 39200 11542 39201
rect 11226 39136 11232 39200
rect 11296 39136 11312 39200
rect 11376 39136 11392 39200
rect 11456 39136 11472 39200
rect 11536 39136 11542 39200
rect 11226 39135 11542 39136
rect 14653 39200 14969 39201
rect 14653 39136 14659 39200
rect 14723 39136 14739 39200
rect 14803 39136 14819 39200
rect 14883 39136 14899 39200
rect 14963 39136 14969 39200
rect 14653 39135 14969 39136
rect 2659 38656 2975 38657
rect 2659 38592 2665 38656
rect 2729 38592 2745 38656
rect 2809 38592 2825 38656
rect 2889 38592 2905 38656
rect 2969 38592 2975 38656
rect 2659 38591 2975 38592
rect 6086 38656 6402 38657
rect 6086 38592 6092 38656
rect 6156 38592 6172 38656
rect 6236 38592 6252 38656
rect 6316 38592 6332 38656
rect 6396 38592 6402 38656
rect 6086 38591 6402 38592
rect 9513 38656 9829 38657
rect 9513 38592 9519 38656
rect 9583 38592 9599 38656
rect 9663 38592 9679 38656
rect 9743 38592 9759 38656
rect 9823 38592 9829 38656
rect 9513 38591 9829 38592
rect 12940 38656 13256 38657
rect 12940 38592 12946 38656
rect 13010 38592 13026 38656
rect 13090 38592 13106 38656
rect 13170 38592 13186 38656
rect 13250 38592 13256 38656
rect 12940 38591 13256 38592
rect 4372 38112 4688 38113
rect 4372 38048 4378 38112
rect 4442 38048 4458 38112
rect 4522 38048 4538 38112
rect 4602 38048 4618 38112
rect 4682 38048 4688 38112
rect 4372 38047 4688 38048
rect 7799 38112 8115 38113
rect 7799 38048 7805 38112
rect 7869 38048 7885 38112
rect 7949 38048 7965 38112
rect 8029 38048 8045 38112
rect 8109 38048 8115 38112
rect 7799 38047 8115 38048
rect 11226 38112 11542 38113
rect 11226 38048 11232 38112
rect 11296 38048 11312 38112
rect 11376 38048 11392 38112
rect 11456 38048 11472 38112
rect 11536 38048 11542 38112
rect 11226 38047 11542 38048
rect 14653 38112 14969 38113
rect 14653 38048 14659 38112
rect 14723 38048 14739 38112
rect 14803 38048 14819 38112
rect 14883 38048 14899 38112
rect 14963 38048 14969 38112
rect 14653 38047 14969 38048
rect 2659 37568 2975 37569
rect 2659 37504 2665 37568
rect 2729 37504 2745 37568
rect 2809 37504 2825 37568
rect 2889 37504 2905 37568
rect 2969 37504 2975 37568
rect 2659 37503 2975 37504
rect 6086 37568 6402 37569
rect 6086 37504 6092 37568
rect 6156 37504 6172 37568
rect 6236 37504 6252 37568
rect 6316 37504 6332 37568
rect 6396 37504 6402 37568
rect 6086 37503 6402 37504
rect 9513 37568 9829 37569
rect 9513 37504 9519 37568
rect 9583 37504 9599 37568
rect 9663 37504 9679 37568
rect 9743 37504 9759 37568
rect 9823 37504 9829 37568
rect 9513 37503 9829 37504
rect 12940 37568 13256 37569
rect 12940 37504 12946 37568
rect 13010 37504 13026 37568
rect 13090 37504 13106 37568
rect 13170 37504 13186 37568
rect 13250 37504 13256 37568
rect 12940 37503 13256 37504
rect 4372 37024 4688 37025
rect 4372 36960 4378 37024
rect 4442 36960 4458 37024
rect 4522 36960 4538 37024
rect 4602 36960 4618 37024
rect 4682 36960 4688 37024
rect 4372 36959 4688 36960
rect 7799 37024 8115 37025
rect 7799 36960 7805 37024
rect 7869 36960 7885 37024
rect 7949 36960 7965 37024
rect 8029 36960 8045 37024
rect 8109 36960 8115 37024
rect 7799 36959 8115 36960
rect 11226 37024 11542 37025
rect 11226 36960 11232 37024
rect 11296 36960 11312 37024
rect 11376 36960 11392 37024
rect 11456 36960 11472 37024
rect 11536 36960 11542 37024
rect 11226 36959 11542 36960
rect 14653 37024 14969 37025
rect 14653 36960 14659 37024
rect 14723 36960 14739 37024
rect 14803 36960 14819 37024
rect 14883 36960 14899 37024
rect 14963 36960 14969 37024
rect 14653 36959 14969 36960
rect 2659 36480 2975 36481
rect 2659 36416 2665 36480
rect 2729 36416 2745 36480
rect 2809 36416 2825 36480
rect 2889 36416 2905 36480
rect 2969 36416 2975 36480
rect 2659 36415 2975 36416
rect 6086 36480 6402 36481
rect 6086 36416 6092 36480
rect 6156 36416 6172 36480
rect 6236 36416 6252 36480
rect 6316 36416 6332 36480
rect 6396 36416 6402 36480
rect 6086 36415 6402 36416
rect 9513 36480 9829 36481
rect 9513 36416 9519 36480
rect 9583 36416 9599 36480
rect 9663 36416 9679 36480
rect 9743 36416 9759 36480
rect 9823 36416 9829 36480
rect 9513 36415 9829 36416
rect 12940 36480 13256 36481
rect 12940 36416 12946 36480
rect 13010 36416 13026 36480
rect 13090 36416 13106 36480
rect 13170 36416 13186 36480
rect 13250 36416 13256 36480
rect 12940 36415 13256 36416
rect 4372 35936 4688 35937
rect 4372 35872 4378 35936
rect 4442 35872 4458 35936
rect 4522 35872 4538 35936
rect 4602 35872 4618 35936
rect 4682 35872 4688 35936
rect 4372 35871 4688 35872
rect 7799 35936 8115 35937
rect 7799 35872 7805 35936
rect 7869 35872 7885 35936
rect 7949 35872 7965 35936
rect 8029 35872 8045 35936
rect 8109 35872 8115 35936
rect 7799 35871 8115 35872
rect 11226 35936 11542 35937
rect 11226 35872 11232 35936
rect 11296 35872 11312 35936
rect 11376 35872 11392 35936
rect 11456 35872 11472 35936
rect 11536 35872 11542 35936
rect 11226 35871 11542 35872
rect 14653 35936 14969 35937
rect 14653 35872 14659 35936
rect 14723 35872 14739 35936
rect 14803 35872 14819 35936
rect 14883 35872 14899 35936
rect 14963 35872 14969 35936
rect 14653 35871 14969 35872
rect 14457 35730 14523 35733
rect 15200 35730 16000 35760
rect 14457 35728 16000 35730
rect 14457 35672 14462 35728
rect 14518 35672 16000 35728
rect 14457 35670 16000 35672
rect 14457 35667 14523 35670
rect 15200 35640 16000 35670
rect 2659 35392 2975 35393
rect 2659 35328 2665 35392
rect 2729 35328 2745 35392
rect 2809 35328 2825 35392
rect 2889 35328 2905 35392
rect 2969 35328 2975 35392
rect 2659 35327 2975 35328
rect 6086 35392 6402 35393
rect 6086 35328 6092 35392
rect 6156 35328 6172 35392
rect 6236 35328 6252 35392
rect 6316 35328 6332 35392
rect 6396 35328 6402 35392
rect 6086 35327 6402 35328
rect 9513 35392 9829 35393
rect 9513 35328 9519 35392
rect 9583 35328 9599 35392
rect 9663 35328 9679 35392
rect 9743 35328 9759 35392
rect 9823 35328 9829 35392
rect 9513 35327 9829 35328
rect 12940 35392 13256 35393
rect 12940 35328 12946 35392
rect 13010 35328 13026 35392
rect 13090 35328 13106 35392
rect 13170 35328 13186 35392
rect 13250 35328 13256 35392
rect 12940 35327 13256 35328
rect 4372 34848 4688 34849
rect 4372 34784 4378 34848
rect 4442 34784 4458 34848
rect 4522 34784 4538 34848
rect 4602 34784 4618 34848
rect 4682 34784 4688 34848
rect 4372 34783 4688 34784
rect 7799 34848 8115 34849
rect 7799 34784 7805 34848
rect 7869 34784 7885 34848
rect 7949 34784 7965 34848
rect 8029 34784 8045 34848
rect 8109 34784 8115 34848
rect 7799 34783 8115 34784
rect 11226 34848 11542 34849
rect 11226 34784 11232 34848
rect 11296 34784 11312 34848
rect 11376 34784 11392 34848
rect 11456 34784 11472 34848
rect 11536 34784 11542 34848
rect 11226 34783 11542 34784
rect 14653 34848 14969 34849
rect 14653 34784 14659 34848
rect 14723 34784 14739 34848
rect 14803 34784 14819 34848
rect 14883 34784 14899 34848
rect 14963 34784 14969 34848
rect 14653 34783 14969 34784
rect 2659 34304 2975 34305
rect 2659 34240 2665 34304
rect 2729 34240 2745 34304
rect 2809 34240 2825 34304
rect 2889 34240 2905 34304
rect 2969 34240 2975 34304
rect 2659 34239 2975 34240
rect 6086 34304 6402 34305
rect 6086 34240 6092 34304
rect 6156 34240 6172 34304
rect 6236 34240 6252 34304
rect 6316 34240 6332 34304
rect 6396 34240 6402 34304
rect 6086 34239 6402 34240
rect 9513 34304 9829 34305
rect 9513 34240 9519 34304
rect 9583 34240 9599 34304
rect 9663 34240 9679 34304
rect 9743 34240 9759 34304
rect 9823 34240 9829 34304
rect 9513 34239 9829 34240
rect 12940 34304 13256 34305
rect 12940 34240 12946 34304
rect 13010 34240 13026 34304
rect 13090 34240 13106 34304
rect 13170 34240 13186 34304
rect 13250 34240 13256 34304
rect 12940 34239 13256 34240
rect 4372 33760 4688 33761
rect 4372 33696 4378 33760
rect 4442 33696 4458 33760
rect 4522 33696 4538 33760
rect 4602 33696 4618 33760
rect 4682 33696 4688 33760
rect 4372 33695 4688 33696
rect 7799 33760 8115 33761
rect 7799 33696 7805 33760
rect 7869 33696 7885 33760
rect 7949 33696 7965 33760
rect 8029 33696 8045 33760
rect 8109 33696 8115 33760
rect 7799 33695 8115 33696
rect 11226 33760 11542 33761
rect 11226 33696 11232 33760
rect 11296 33696 11312 33760
rect 11376 33696 11392 33760
rect 11456 33696 11472 33760
rect 11536 33696 11542 33760
rect 11226 33695 11542 33696
rect 14653 33760 14969 33761
rect 14653 33696 14659 33760
rect 14723 33696 14739 33760
rect 14803 33696 14819 33760
rect 14883 33696 14899 33760
rect 14963 33696 14969 33760
rect 14653 33695 14969 33696
rect 2659 33216 2975 33217
rect 2659 33152 2665 33216
rect 2729 33152 2745 33216
rect 2809 33152 2825 33216
rect 2889 33152 2905 33216
rect 2969 33152 2975 33216
rect 2659 33151 2975 33152
rect 6086 33216 6402 33217
rect 6086 33152 6092 33216
rect 6156 33152 6172 33216
rect 6236 33152 6252 33216
rect 6316 33152 6332 33216
rect 6396 33152 6402 33216
rect 6086 33151 6402 33152
rect 9513 33216 9829 33217
rect 9513 33152 9519 33216
rect 9583 33152 9599 33216
rect 9663 33152 9679 33216
rect 9743 33152 9759 33216
rect 9823 33152 9829 33216
rect 9513 33151 9829 33152
rect 12940 33216 13256 33217
rect 12940 33152 12946 33216
rect 13010 33152 13026 33216
rect 13090 33152 13106 33216
rect 13170 33152 13186 33216
rect 13250 33152 13256 33216
rect 12940 33151 13256 33152
rect 4372 32672 4688 32673
rect 4372 32608 4378 32672
rect 4442 32608 4458 32672
rect 4522 32608 4538 32672
rect 4602 32608 4618 32672
rect 4682 32608 4688 32672
rect 4372 32607 4688 32608
rect 7799 32672 8115 32673
rect 7799 32608 7805 32672
rect 7869 32608 7885 32672
rect 7949 32608 7965 32672
rect 8029 32608 8045 32672
rect 8109 32608 8115 32672
rect 7799 32607 8115 32608
rect 11226 32672 11542 32673
rect 11226 32608 11232 32672
rect 11296 32608 11312 32672
rect 11376 32608 11392 32672
rect 11456 32608 11472 32672
rect 11536 32608 11542 32672
rect 11226 32607 11542 32608
rect 14653 32672 14969 32673
rect 14653 32608 14659 32672
rect 14723 32608 14739 32672
rect 14803 32608 14819 32672
rect 14883 32608 14899 32672
rect 14963 32608 14969 32672
rect 14653 32607 14969 32608
rect 2659 32128 2975 32129
rect 2659 32064 2665 32128
rect 2729 32064 2745 32128
rect 2809 32064 2825 32128
rect 2889 32064 2905 32128
rect 2969 32064 2975 32128
rect 2659 32063 2975 32064
rect 6086 32128 6402 32129
rect 6086 32064 6092 32128
rect 6156 32064 6172 32128
rect 6236 32064 6252 32128
rect 6316 32064 6332 32128
rect 6396 32064 6402 32128
rect 6086 32063 6402 32064
rect 9513 32128 9829 32129
rect 9513 32064 9519 32128
rect 9583 32064 9599 32128
rect 9663 32064 9679 32128
rect 9743 32064 9759 32128
rect 9823 32064 9829 32128
rect 9513 32063 9829 32064
rect 12940 32128 13256 32129
rect 12940 32064 12946 32128
rect 13010 32064 13026 32128
rect 13090 32064 13106 32128
rect 13170 32064 13186 32128
rect 13250 32064 13256 32128
rect 12940 32063 13256 32064
rect 4372 31584 4688 31585
rect 4372 31520 4378 31584
rect 4442 31520 4458 31584
rect 4522 31520 4538 31584
rect 4602 31520 4618 31584
rect 4682 31520 4688 31584
rect 4372 31519 4688 31520
rect 7799 31584 8115 31585
rect 7799 31520 7805 31584
rect 7869 31520 7885 31584
rect 7949 31520 7965 31584
rect 8029 31520 8045 31584
rect 8109 31520 8115 31584
rect 7799 31519 8115 31520
rect 11226 31584 11542 31585
rect 11226 31520 11232 31584
rect 11296 31520 11312 31584
rect 11376 31520 11392 31584
rect 11456 31520 11472 31584
rect 11536 31520 11542 31584
rect 11226 31519 11542 31520
rect 14653 31584 14969 31585
rect 14653 31520 14659 31584
rect 14723 31520 14739 31584
rect 14803 31520 14819 31584
rect 14883 31520 14899 31584
rect 14963 31520 14969 31584
rect 14653 31519 14969 31520
rect 2659 31040 2975 31041
rect 2659 30976 2665 31040
rect 2729 30976 2745 31040
rect 2809 30976 2825 31040
rect 2889 30976 2905 31040
rect 2969 30976 2975 31040
rect 2659 30975 2975 30976
rect 6086 31040 6402 31041
rect 6086 30976 6092 31040
rect 6156 30976 6172 31040
rect 6236 30976 6252 31040
rect 6316 30976 6332 31040
rect 6396 30976 6402 31040
rect 6086 30975 6402 30976
rect 9513 31040 9829 31041
rect 9513 30976 9519 31040
rect 9583 30976 9599 31040
rect 9663 30976 9679 31040
rect 9743 30976 9759 31040
rect 9823 30976 9829 31040
rect 9513 30975 9829 30976
rect 12940 31040 13256 31041
rect 12940 30976 12946 31040
rect 13010 30976 13026 31040
rect 13090 30976 13106 31040
rect 13170 30976 13186 31040
rect 13250 30976 13256 31040
rect 12940 30975 13256 30976
rect 4372 30496 4688 30497
rect 4372 30432 4378 30496
rect 4442 30432 4458 30496
rect 4522 30432 4538 30496
rect 4602 30432 4618 30496
rect 4682 30432 4688 30496
rect 4372 30431 4688 30432
rect 7799 30496 8115 30497
rect 7799 30432 7805 30496
rect 7869 30432 7885 30496
rect 7949 30432 7965 30496
rect 8029 30432 8045 30496
rect 8109 30432 8115 30496
rect 7799 30431 8115 30432
rect 11226 30496 11542 30497
rect 11226 30432 11232 30496
rect 11296 30432 11312 30496
rect 11376 30432 11392 30496
rect 11456 30432 11472 30496
rect 11536 30432 11542 30496
rect 11226 30431 11542 30432
rect 14653 30496 14969 30497
rect 14653 30432 14659 30496
rect 14723 30432 14739 30496
rect 14803 30432 14819 30496
rect 14883 30432 14899 30496
rect 14963 30432 14969 30496
rect 14653 30431 14969 30432
rect 2659 29952 2975 29953
rect 2659 29888 2665 29952
rect 2729 29888 2745 29952
rect 2809 29888 2825 29952
rect 2889 29888 2905 29952
rect 2969 29888 2975 29952
rect 2659 29887 2975 29888
rect 6086 29952 6402 29953
rect 6086 29888 6092 29952
rect 6156 29888 6172 29952
rect 6236 29888 6252 29952
rect 6316 29888 6332 29952
rect 6396 29888 6402 29952
rect 6086 29887 6402 29888
rect 9513 29952 9829 29953
rect 9513 29888 9519 29952
rect 9583 29888 9599 29952
rect 9663 29888 9679 29952
rect 9743 29888 9759 29952
rect 9823 29888 9829 29952
rect 9513 29887 9829 29888
rect 12940 29952 13256 29953
rect 12940 29888 12946 29952
rect 13010 29888 13026 29952
rect 13090 29888 13106 29952
rect 13170 29888 13186 29952
rect 13250 29888 13256 29952
rect 12940 29887 13256 29888
rect 4372 29408 4688 29409
rect 4372 29344 4378 29408
rect 4442 29344 4458 29408
rect 4522 29344 4538 29408
rect 4602 29344 4618 29408
rect 4682 29344 4688 29408
rect 4372 29343 4688 29344
rect 7799 29408 8115 29409
rect 7799 29344 7805 29408
rect 7869 29344 7885 29408
rect 7949 29344 7965 29408
rect 8029 29344 8045 29408
rect 8109 29344 8115 29408
rect 7799 29343 8115 29344
rect 11226 29408 11542 29409
rect 11226 29344 11232 29408
rect 11296 29344 11312 29408
rect 11376 29344 11392 29408
rect 11456 29344 11472 29408
rect 11536 29344 11542 29408
rect 11226 29343 11542 29344
rect 14653 29408 14969 29409
rect 14653 29344 14659 29408
rect 14723 29344 14739 29408
rect 14803 29344 14819 29408
rect 14883 29344 14899 29408
rect 14963 29344 14969 29408
rect 14653 29343 14969 29344
rect 2659 28864 2975 28865
rect 2659 28800 2665 28864
rect 2729 28800 2745 28864
rect 2809 28800 2825 28864
rect 2889 28800 2905 28864
rect 2969 28800 2975 28864
rect 2659 28799 2975 28800
rect 6086 28864 6402 28865
rect 6086 28800 6092 28864
rect 6156 28800 6172 28864
rect 6236 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6402 28864
rect 6086 28799 6402 28800
rect 9513 28864 9829 28865
rect 9513 28800 9519 28864
rect 9583 28800 9599 28864
rect 9663 28800 9679 28864
rect 9743 28800 9759 28864
rect 9823 28800 9829 28864
rect 9513 28799 9829 28800
rect 12940 28864 13256 28865
rect 12940 28800 12946 28864
rect 13010 28800 13026 28864
rect 13090 28800 13106 28864
rect 13170 28800 13186 28864
rect 13250 28800 13256 28864
rect 12940 28799 13256 28800
rect 4372 28320 4688 28321
rect 4372 28256 4378 28320
rect 4442 28256 4458 28320
rect 4522 28256 4538 28320
rect 4602 28256 4618 28320
rect 4682 28256 4688 28320
rect 4372 28255 4688 28256
rect 7799 28320 8115 28321
rect 7799 28256 7805 28320
rect 7869 28256 7885 28320
rect 7949 28256 7965 28320
rect 8029 28256 8045 28320
rect 8109 28256 8115 28320
rect 7799 28255 8115 28256
rect 11226 28320 11542 28321
rect 11226 28256 11232 28320
rect 11296 28256 11312 28320
rect 11376 28256 11392 28320
rect 11456 28256 11472 28320
rect 11536 28256 11542 28320
rect 11226 28255 11542 28256
rect 14653 28320 14969 28321
rect 14653 28256 14659 28320
rect 14723 28256 14739 28320
rect 14803 28256 14819 28320
rect 14883 28256 14899 28320
rect 14963 28256 14969 28320
rect 14653 28255 14969 28256
rect 14457 27842 14523 27845
rect 15200 27842 16000 27872
rect 14457 27840 16000 27842
rect 14457 27784 14462 27840
rect 14518 27784 16000 27840
rect 14457 27782 16000 27784
rect 14457 27779 14523 27782
rect 2659 27776 2975 27777
rect 2659 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2975 27776
rect 2659 27711 2975 27712
rect 6086 27776 6402 27777
rect 6086 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6402 27776
rect 6086 27711 6402 27712
rect 9513 27776 9829 27777
rect 9513 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9829 27776
rect 9513 27711 9829 27712
rect 12940 27776 13256 27777
rect 12940 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13256 27776
rect 15200 27752 16000 27782
rect 12940 27711 13256 27712
rect 4372 27232 4688 27233
rect 4372 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4688 27232
rect 4372 27167 4688 27168
rect 7799 27232 8115 27233
rect 7799 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8115 27232
rect 7799 27167 8115 27168
rect 11226 27232 11542 27233
rect 11226 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11542 27232
rect 11226 27167 11542 27168
rect 14653 27232 14969 27233
rect 14653 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14969 27232
rect 14653 27167 14969 27168
rect 2659 26688 2975 26689
rect 2659 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2975 26688
rect 2659 26623 2975 26624
rect 6086 26688 6402 26689
rect 6086 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6402 26688
rect 6086 26623 6402 26624
rect 9513 26688 9829 26689
rect 9513 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9829 26688
rect 9513 26623 9829 26624
rect 12940 26688 13256 26689
rect 12940 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13256 26688
rect 12940 26623 13256 26624
rect 4372 26144 4688 26145
rect 4372 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4688 26144
rect 4372 26079 4688 26080
rect 7799 26144 8115 26145
rect 7799 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8115 26144
rect 7799 26079 8115 26080
rect 11226 26144 11542 26145
rect 11226 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11542 26144
rect 11226 26079 11542 26080
rect 14653 26144 14969 26145
rect 14653 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14969 26144
rect 14653 26079 14969 26080
rect 2659 25600 2975 25601
rect 2659 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2975 25600
rect 2659 25535 2975 25536
rect 6086 25600 6402 25601
rect 6086 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6402 25600
rect 6086 25535 6402 25536
rect 9513 25600 9829 25601
rect 9513 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9829 25600
rect 9513 25535 9829 25536
rect 12940 25600 13256 25601
rect 12940 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13256 25600
rect 12940 25535 13256 25536
rect 4372 25056 4688 25057
rect 4372 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4688 25056
rect 4372 24991 4688 24992
rect 7799 25056 8115 25057
rect 7799 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8115 25056
rect 7799 24991 8115 24992
rect 11226 25056 11542 25057
rect 11226 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11542 25056
rect 11226 24991 11542 24992
rect 14653 25056 14969 25057
rect 14653 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14969 25056
rect 14653 24991 14969 24992
rect 2659 24512 2975 24513
rect 2659 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2975 24512
rect 2659 24447 2975 24448
rect 6086 24512 6402 24513
rect 6086 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6402 24512
rect 6086 24447 6402 24448
rect 9513 24512 9829 24513
rect 9513 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9829 24512
rect 9513 24447 9829 24448
rect 12940 24512 13256 24513
rect 12940 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13256 24512
rect 12940 24447 13256 24448
rect 4372 23968 4688 23969
rect 4372 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4688 23968
rect 4372 23903 4688 23904
rect 7799 23968 8115 23969
rect 7799 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8115 23968
rect 7799 23903 8115 23904
rect 11226 23968 11542 23969
rect 11226 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11542 23968
rect 11226 23903 11542 23904
rect 14653 23968 14969 23969
rect 14653 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14969 23968
rect 14653 23903 14969 23904
rect 2659 23424 2975 23425
rect 2659 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2975 23424
rect 2659 23359 2975 23360
rect 6086 23424 6402 23425
rect 6086 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6402 23424
rect 6086 23359 6402 23360
rect 9513 23424 9829 23425
rect 9513 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9829 23424
rect 9513 23359 9829 23360
rect 12940 23424 13256 23425
rect 12940 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13256 23424
rect 12940 23359 13256 23360
rect 4372 22880 4688 22881
rect 4372 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4688 22880
rect 4372 22815 4688 22816
rect 7799 22880 8115 22881
rect 7799 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8115 22880
rect 7799 22815 8115 22816
rect 11226 22880 11542 22881
rect 11226 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11542 22880
rect 11226 22815 11542 22816
rect 14653 22880 14969 22881
rect 14653 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14969 22880
rect 14653 22815 14969 22816
rect 2659 22336 2975 22337
rect 2659 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2975 22336
rect 2659 22271 2975 22272
rect 6086 22336 6402 22337
rect 6086 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6402 22336
rect 6086 22271 6402 22272
rect 9513 22336 9829 22337
rect 9513 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9829 22336
rect 9513 22271 9829 22272
rect 12940 22336 13256 22337
rect 12940 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13256 22336
rect 12940 22271 13256 22272
rect 4372 21792 4688 21793
rect 4372 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4688 21792
rect 4372 21727 4688 21728
rect 7799 21792 8115 21793
rect 7799 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8115 21792
rect 7799 21727 8115 21728
rect 11226 21792 11542 21793
rect 11226 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11542 21792
rect 11226 21727 11542 21728
rect 14653 21792 14969 21793
rect 14653 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14969 21792
rect 14653 21727 14969 21728
rect 2659 21248 2975 21249
rect 2659 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2975 21248
rect 2659 21183 2975 21184
rect 6086 21248 6402 21249
rect 6086 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6402 21248
rect 6086 21183 6402 21184
rect 9513 21248 9829 21249
rect 9513 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9829 21248
rect 9513 21183 9829 21184
rect 12940 21248 13256 21249
rect 12940 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13256 21248
rect 12940 21183 13256 21184
rect 4372 20704 4688 20705
rect 4372 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4688 20704
rect 4372 20639 4688 20640
rect 7799 20704 8115 20705
rect 7799 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8115 20704
rect 7799 20639 8115 20640
rect 11226 20704 11542 20705
rect 11226 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11542 20704
rect 11226 20639 11542 20640
rect 14653 20704 14969 20705
rect 14653 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14969 20704
rect 14653 20639 14969 20640
rect 2659 20160 2975 20161
rect 2659 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2975 20160
rect 2659 20095 2975 20096
rect 6086 20160 6402 20161
rect 6086 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6402 20160
rect 6086 20095 6402 20096
rect 9513 20160 9829 20161
rect 9513 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9829 20160
rect 9513 20095 9829 20096
rect 12940 20160 13256 20161
rect 12940 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13256 20160
rect 12940 20095 13256 20096
rect 14457 19954 14523 19957
rect 15200 19954 16000 19984
rect 14457 19952 16000 19954
rect 14457 19896 14462 19952
rect 14518 19896 16000 19952
rect 14457 19894 16000 19896
rect 14457 19891 14523 19894
rect 15200 19864 16000 19894
rect 4372 19616 4688 19617
rect 4372 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4688 19616
rect 4372 19551 4688 19552
rect 7799 19616 8115 19617
rect 7799 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8115 19616
rect 7799 19551 8115 19552
rect 11226 19616 11542 19617
rect 11226 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11542 19616
rect 11226 19551 11542 19552
rect 14653 19616 14969 19617
rect 14653 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14969 19616
rect 14653 19551 14969 19552
rect 2659 19072 2975 19073
rect 2659 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2975 19072
rect 2659 19007 2975 19008
rect 6086 19072 6402 19073
rect 6086 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6402 19072
rect 6086 19007 6402 19008
rect 9513 19072 9829 19073
rect 9513 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9829 19072
rect 9513 19007 9829 19008
rect 12940 19072 13256 19073
rect 12940 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13256 19072
rect 12940 19007 13256 19008
rect 4372 18528 4688 18529
rect 4372 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4688 18528
rect 4372 18463 4688 18464
rect 7799 18528 8115 18529
rect 7799 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8115 18528
rect 7799 18463 8115 18464
rect 11226 18528 11542 18529
rect 11226 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11542 18528
rect 11226 18463 11542 18464
rect 14653 18528 14969 18529
rect 14653 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14969 18528
rect 14653 18463 14969 18464
rect 2659 17984 2975 17985
rect 2659 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2975 17984
rect 2659 17919 2975 17920
rect 6086 17984 6402 17985
rect 6086 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6402 17984
rect 6086 17919 6402 17920
rect 9513 17984 9829 17985
rect 9513 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9829 17984
rect 9513 17919 9829 17920
rect 12940 17984 13256 17985
rect 12940 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13256 17984
rect 12940 17919 13256 17920
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 12940 16831 13256 16832
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 14653 16287 14969 16288
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 14653 15199 14969 15200
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 14457 12202 14523 12205
rect 14457 12200 15210 12202
rect 14457 12144 14462 12200
rect 14518 12144 15210 12200
rect 14457 12142 15210 12144
rect 14457 12139 14523 12142
rect 15150 12096 15210 12142
rect 15150 12006 16000 12096
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 15200 11976 16000 12006
rect 14653 11935 14969 11936
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 12940 10303 13256 10304
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 14653 9759 14969 9760
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 14653 8671 14969 8672
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 12940 7039 13256 7040
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 14457 4178 14523 4181
rect 15200 4178 16000 4208
rect 14457 4176 16000 4178
rect 14457 4120 14462 4176
rect 14518 4120 16000 4176
rect 14457 4118 16000 4120
rect 14457 4115 14523 4118
rect 15200 4088 16000 4118
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
<< via3 >>
rect 4378 45724 4442 45728
rect 4378 45668 4382 45724
rect 4382 45668 4438 45724
rect 4438 45668 4442 45724
rect 4378 45664 4442 45668
rect 4458 45724 4522 45728
rect 4458 45668 4462 45724
rect 4462 45668 4518 45724
rect 4518 45668 4522 45724
rect 4458 45664 4522 45668
rect 4538 45724 4602 45728
rect 4538 45668 4542 45724
rect 4542 45668 4598 45724
rect 4598 45668 4602 45724
rect 4538 45664 4602 45668
rect 4618 45724 4682 45728
rect 4618 45668 4622 45724
rect 4622 45668 4678 45724
rect 4678 45668 4682 45724
rect 4618 45664 4682 45668
rect 7805 45724 7869 45728
rect 7805 45668 7809 45724
rect 7809 45668 7865 45724
rect 7865 45668 7869 45724
rect 7805 45664 7869 45668
rect 7885 45724 7949 45728
rect 7885 45668 7889 45724
rect 7889 45668 7945 45724
rect 7945 45668 7949 45724
rect 7885 45664 7949 45668
rect 7965 45724 8029 45728
rect 7965 45668 7969 45724
rect 7969 45668 8025 45724
rect 8025 45668 8029 45724
rect 7965 45664 8029 45668
rect 8045 45724 8109 45728
rect 8045 45668 8049 45724
rect 8049 45668 8105 45724
rect 8105 45668 8109 45724
rect 8045 45664 8109 45668
rect 11232 45724 11296 45728
rect 11232 45668 11236 45724
rect 11236 45668 11292 45724
rect 11292 45668 11296 45724
rect 11232 45664 11296 45668
rect 11312 45724 11376 45728
rect 11312 45668 11316 45724
rect 11316 45668 11372 45724
rect 11372 45668 11376 45724
rect 11312 45664 11376 45668
rect 11392 45724 11456 45728
rect 11392 45668 11396 45724
rect 11396 45668 11452 45724
rect 11452 45668 11456 45724
rect 11392 45664 11456 45668
rect 11472 45724 11536 45728
rect 11472 45668 11476 45724
rect 11476 45668 11532 45724
rect 11532 45668 11536 45724
rect 11472 45664 11536 45668
rect 14659 45724 14723 45728
rect 14659 45668 14663 45724
rect 14663 45668 14719 45724
rect 14719 45668 14723 45724
rect 14659 45664 14723 45668
rect 14739 45724 14803 45728
rect 14739 45668 14743 45724
rect 14743 45668 14799 45724
rect 14799 45668 14803 45724
rect 14739 45664 14803 45668
rect 14819 45724 14883 45728
rect 14819 45668 14823 45724
rect 14823 45668 14879 45724
rect 14879 45668 14883 45724
rect 14819 45664 14883 45668
rect 14899 45724 14963 45728
rect 14899 45668 14903 45724
rect 14903 45668 14959 45724
rect 14959 45668 14963 45724
rect 14899 45664 14963 45668
rect 2665 45180 2729 45184
rect 2665 45124 2669 45180
rect 2669 45124 2725 45180
rect 2725 45124 2729 45180
rect 2665 45120 2729 45124
rect 2745 45180 2809 45184
rect 2745 45124 2749 45180
rect 2749 45124 2805 45180
rect 2805 45124 2809 45180
rect 2745 45120 2809 45124
rect 2825 45180 2889 45184
rect 2825 45124 2829 45180
rect 2829 45124 2885 45180
rect 2885 45124 2889 45180
rect 2825 45120 2889 45124
rect 2905 45180 2969 45184
rect 2905 45124 2909 45180
rect 2909 45124 2965 45180
rect 2965 45124 2969 45180
rect 2905 45120 2969 45124
rect 6092 45180 6156 45184
rect 6092 45124 6096 45180
rect 6096 45124 6152 45180
rect 6152 45124 6156 45180
rect 6092 45120 6156 45124
rect 6172 45180 6236 45184
rect 6172 45124 6176 45180
rect 6176 45124 6232 45180
rect 6232 45124 6236 45180
rect 6172 45120 6236 45124
rect 6252 45180 6316 45184
rect 6252 45124 6256 45180
rect 6256 45124 6312 45180
rect 6312 45124 6316 45180
rect 6252 45120 6316 45124
rect 6332 45180 6396 45184
rect 6332 45124 6336 45180
rect 6336 45124 6392 45180
rect 6392 45124 6396 45180
rect 6332 45120 6396 45124
rect 9519 45180 9583 45184
rect 9519 45124 9523 45180
rect 9523 45124 9579 45180
rect 9579 45124 9583 45180
rect 9519 45120 9583 45124
rect 9599 45180 9663 45184
rect 9599 45124 9603 45180
rect 9603 45124 9659 45180
rect 9659 45124 9663 45180
rect 9599 45120 9663 45124
rect 9679 45180 9743 45184
rect 9679 45124 9683 45180
rect 9683 45124 9739 45180
rect 9739 45124 9743 45180
rect 9679 45120 9743 45124
rect 9759 45180 9823 45184
rect 9759 45124 9763 45180
rect 9763 45124 9819 45180
rect 9819 45124 9823 45180
rect 9759 45120 9823 45124
rect 12946 45180 13010 45184
rect 12946 45124 12950 45180
rect 12950 45124 13006 45180
rect 13006 45124 13010 45180
rect 12946 45120 13010 45124
rect 13026 45180 13090 45184
rect 13026 45124 13030 45180
rect 13030 45124 13086 45180
rect 13086 45124 13090 45180
rect 13026 45120 13090 45124
rect 13106 45180 13170 45184
rect 13106 45124 13110 45180
rect 13110 45124 13166 45180
rect 13166 45124 13170 45180
rect 13106 45120 13170 45124
rect 13186 45180 13250 45184
rect 13186 45124 13190 45180
rect 13190 45124 13246 45180
rect 13246 45124 13250 45180
rect 13186 45120 13250 45124
rect 4378 44636 4442 44640
rect 4378 44580 4382 44636
rect 4382 44580 4438 44636
rect 4438 44580 4442 44636
rect 4378 44576 4442 44580
rect 4458 44636 4522 44640
rect 4458 44580 4462 44636
rect 4462 44580 4518 44636
rect 4518 44580 4522 44636
rect 4458 44576 4522 44580
rect 4538 44636 4602 44640
rect 4538 44580 4542 44636
rect 4542 44580 4598 44636
rect 4598 44580 4602 44636
rect 4538 44576 4602 44580
rect 4618 44636 4682 44640
rect 4618 44580 4622 44636
rect 4622 44580 4678 44636
rect 4678 44580 4682 44636
rect 4618 44576 4682 44580
rect 7805 44636 7869 44640
rect 7805 44580 7809 44636
rect 7809 44580 7865 44636
rect 7865 44580 7869 44636
rect 7805 44576 7869 44580
rect 7885 44636 7949 44640
rect 7885 44580 7889 44636
rect 7889 44580 7945 44636
rect 7945 44580 7949 44636
rect 7885 44576 7949 44580
rect 7965 44636 8029 44640
rect 7965 44580 7969 44636
rect 7969 44580 8025 44636
rect 8025 44580 8029 44636
rect 7965 44576 8029 44580
rect 8045 44636 8109 44640
rect 8045 44580 8049 44636
rect 8049 44580 8105 44636
rect 8105 44580 8109 44636
rect 8045 44576 8109 44580
rect 11232 44636 11296 44640
rect 11232 44580 11236 44636
rect 11236 44580 11292 44636
rect 11292 44580 11296 44636
rect 11232 44576 11296 44580
rect 11312 44636 11376 44640
rect 11312 44580 11316 44636
rect 11316 44580 11372 44636
rect 11372 44580 11376 44636
rect 11312 44576 11376 44580
rect 11392 44636 11456 44640
rect 11392 44580 11396 44636
rect 11396 44580 11452 44636
rect 11452 44580 11456 44636
rect 11392 44576 11456 44580
rect 11472 44636 11536 44640
rect 11472 44580 11476 44636
rect 11476 44580 11532 44636
rect 11532 44580 11536 44636
rect 11472 44576 11536 44580
rect 14659 44636 14723 44640
rect 14659 44580 14663 44636
rect 14663 44580 14719 44636
rect 14719 44580 14723 44636
rect 14659 44576 14723 44580
rect 14739 44636 14803 44640
rect 14739 44580 14743 44636
rect 14743 44580 14799 44636
rect 14799 44580 14803 44636
rect 14739 44576 14803 44580
rect 14819 44636 14883 44640
rect 14819 44580 14823 44636
rect 14823 44580 14879 44636
rect 14879 44580 14883 44636
rect 14819 44576 14883 44580
rect 14899 44636 14963 44640
rect 14899 44580 14903 44636
rect 14903 44580 14959 44636
rect 14959 44580 14963 44636
rect 14899 44576 14963 44580
rect 2665 44092 2729 44096
rect 2665 44036 2669 44092
rect 2669 44036 2725 44092
rect 2725 44036 2729 44092
rect 2665 44032 2729 44036
rect 2745 44092 2809 44096
rect 2745 44036 2749 44092
rect 2749 44036 2805 44092
rect 2805 44036 2809 44092
rect 2745 44032 2809 44036
rect 2825 44092 2889 44096
rect 2825 44036 2829 44092
rect 2829 44036 2885 44092
rect 2885 44036 2889 44092
rect 2825 44032 2889 44036
rect 2905 44092 2969 44096
rect 2905 44036 2909 44092
rect 2909 44036 2965 44092
rect 2965 44036 2969 44092
rect 2905 44032 2969 44036
rect 6092 44092 6156 44096
rect 6092 44036 6096 44092
rect 6096 44036 6152 44092
rect 6152 44036 6156 44092
rect 6092 44032 6156 44036
rect 6172 44092 6236 44096
rect 6172 44036 6176 44092
rect 6176 44036 6232 44092
rect 6232 44036 6236 44092
rect 6172 44032 6236 44036
rect 6252 44092 6316 44096
rect 6252 44036 6256 44092
rect 6256 44036 6312 44092
rect 6312 44036 6316 44092
rect 6252 44032 6316 44036
rect 6332 44092 6396 44096
rect 6332 44036 6336 44092
rect 6336 44036 6392 44092
rect 6392 44036 6396 44092
rect 6332 44032 6396 44036
rect 9519 44092 9583 44096
rect 9519 44036 9523 44092
rect 9523 44036 9579 44092
rect 9579 44036 9583 44092
rect 9519 44032 9583 44036
rect 9599 44092 9663 44096
rect 9599 44036 9603 44092
rect 9603 44036 9659 44092
rect 9659 44036 9663 44092
rect 9599 44032 9663 44036
rect 9679 44092 9743 44096
rect 9679 44036 9683 44092
rect 9683 44036 9739 44092
rect 9739 44036 9743 44092
rect 9679 44032 9743 44036
rect 9759 44092 9823 44096
rect 9759 44036 9763 44092
rect 9763 44036 9819 44092
rect 9819 44036 9823 44092
rect 9759 44032 9823 44036
rect 12946 44092 13010 44096
rect 12946 44036 12950 44092
rect 12950 44036 13006 44092
rect 13006 44036 13010 44092
rect 12946 44032 13010 44036
rect 13026 44092 13090 44096
rect 13026 44036 13030 44092
rect 13030 44036 13086 44092
rect 13086 44036 13090 44092
rect 13026 44032 13090 44036
rect 13106 44092 13170 44096
rect 13106 44036 13110 44092
rect 13110 44036 13166 44092
rect 13166 44036 13170 44092
rect 13106 44032 13170 44036
rect 13186 44092 13250 44096
rect 13186 44036 13190 44092
rect 13190 44036 13246 44092
rect 13246 44036 13250 44092
rect 13186 44032 13250 44036
rect 4378 43548 4442 43552
rect 4378 43492 4382 43548
rect 4382 43492 4438 43548
rect 4438 43492 4442 43548
rect 4378 43488 4442 43492
rect 4458 43548 4522 43552
rect 4458 43492 4462 43548
rect 4462 43492 4518 43548
rect 4518 43492 4522 43548
rect 4458 43488 4522 43492
rect 4538 43548 4602 43552
rect 4538 43492 4542 43548
rect 4542 43492 4598 43548
rect 4598 43492 4602 43548
rect 4538 43488 4602 43492
rect 4618 43548 4682 43552
rect 4618 43492 4622 43548
rect 4622 43492 4678 43548
rect 4678 43492 4682 43548
rect 4618 43488 4682 43492
rect 7805 43548 7869 43552
rect 7805 43492 7809 43548
rect 7809 43492 7865 43548
rect 7865 43492 7869 43548
rect 7805 43488 7869 43492
rect 7885 43548 7949 43552
rect 7885 43492 7889 43548
rect 7889 43492 7945 43548
rect 7945 43492 7949 43548
rect 7885 43488 7949 43492
rect 7965 43548 8029 43552
rect 7965 43492 7969 43548
rect 7969 43492 8025 43548
rect 8025 43492 8029 43548
rect 7965 43488 8029 43492
rect 8045 43548 8109 43552
rect 8045 43492 8049 43548
rect 8049 43492 8105 43548
rect 8105 43492 8109 43548
rect 8045 43488 8109 43492
rect 11232 43548 11296 43552
rect 11232 43492 11236 43548
rect 11236 43492 11292 43548
rect 11292 43492 11296 43548
rect 11232 43488 11296 43492
rect 11312 43548 11376 43552
rect 11312 43492 11316 43548
rect 11316 43492 11372 43548
rect 11372 43492 11376 43548
rect 11312 43488 11376 43492
rect 11392 43548 11456 43552
rect 11392 43492 11396 43548
rect 11396 43492 11452 43548
rect 11452 43492 11456 43548
rect 11392 43488 11456 43492
rect 11472 43548 11536 43552
rect 11472 43492 11476 43548
rect 11476 43492 11532 43548
rect 11532 43492 11536 43548
rect 11472 43488 11536 43492
rect 14659 43548 14723 43552
rect 14659 43492 14663 43548
rect 14663 43492 14719 43548
rect 14719 43492 14723 43548
rect 14659 43488 14723 43492
rect 14739 43548 14803 43552
rect 14739 43492 14743 43548
rect 14743 43492 14799 43548
rect 14799 43492 14803 43548
rect 14739 43488 14803 43492
rect 14819 43548 14883 43552
rect 14819 43492 14823 43548
rect 14823 43492 14879 43548
rect 14879 43492 14883 43548
rect 14819 43488 14883 43492
rect 14899 43548 14963 43552
rect 14899 43492 14903 43548
rect 14903 43492 14959 43548
rect 14959 43492 14963 43548
rect 14899 43488 14963 43492
rect 2665 43004 2729 43008
rect 2665 42948 2669 43004
rect 2669 42948 2725 43004
rect 2725 42948 2729 43004
rect 2665 42944 2729 42948
rect 2745 43004 2809 43008
rect 2745 42948 2749 43004
rect 2749 42948 2805 43004
rect 2805 42948 2809 43004
rect 2745 42944 2809 42948
rect 2825 43004 2889 43008
rect 2825 42948 2829 43004
rect 2829 42948 2885 43004
rect 2885 42948 2889 43004
rect 2825 42944 2889 42948
rect 2905 43004 2969 43008
rect 2905 42948 2909 43004
rect 2909 42948 2965 43004
rect 2965 42948 2969 43004
rect 2905 42944 2969 42948
rect 6092 43004 6156 43008
rect 6092 42948 6096 43004
rect 6096 42948 6152 43004
rect 6152 42948 6156 43004
rect 6092 42944 6156 42948
rect 6172 43004 6236 43008
rect 6172 42948 6176 43004
rect 6176 42948 6232 43004
rect 6232 42948 6236 43004
rect 6172 42944 6236 42948
rect 6252 43004 6316 43008
rect 6252 42948 6256 43004
rect 6256 42948 6312 43004
rect 6312 42948 6316 43004
rect 6252 42944 6316 42948
rect 6332 43004 6396 43008
rect 6332 42948 6336 43004
rect 6336 42948 6392 43004
rect 6392 42948 6396 43004
rect 6332 42944 6396 42948
rect 9519 43004 9583 43008
rect 9519 42948 9523 43004
rect 9523 42948 9579 43004
rect 9579 42948 9583 43004
rect 9519 42944 9583 42948
rect 9599 43004 9663 43008
rect 9599 42948 9603 43004
rect 9603 42948 9659 43004
rect 9659 42948 9663 43004
rect 9599 42944 9663 42948
rect 9679 43004 9743 43008
rect 9679 42948 9683 43004
rect 9683 42948 9739 43004
rect 9739 42948 9743 43004
rect 9679 42944 9743 42948
rect 9759 43004 9823 43008
rect 9759 42948 9763 43004
rect 9763 42948 9819 43004
rect 9819 42948 9823 43004
rect 9759 42944 9823 42948
rect 12946 43004 13010 43008
rect 12946 42948 12950 43004
rect 12950 42948 13006 43004
rect 13006 42948 13010 43004
rect 12946 42944 13010 42948
rect 13026 43004 13090 43008
rect 13026 42948 13030 43004
rect 13030 42948 13086 43004
rect 13086 42948 13090 43004
rect 13026 42944 13090 42948
rect 13106 43004 13170 43008
rect 13106 42948 13110 43004
rect 13110 42948 13166 43004
rect 13166 42948 13170 43004
rect 13106 42944 13170 42948
rect 13186 43004 13250 43008
rect 13186 42948 13190 43004
rect 13190 42948 13246 43004
rect 13246 42948 13250 43004
rect 13186 42944 13250 42948
rect 4378 42460 4442 42464
rect 4378 42404 4382 42460
rect 4382 42404 4438 42460
rect 4438 42404 4442 42460
rect 4378 42400 4442 42404
rect 4458 42460 4522 42464
rect 4458 42404 4462 42460
rect 4462 42404 4518 42460
rect 4518 42404 4522 42460
rect 4458 42400 4522 42404
rect 4538 42460 4602 42464
rect 4538 42404 4542 42460
rect 4542 42404 4598 42460
rect 4598 42404 4602 42460
rect 4538 42400 4602 42404
rect 4618 42460 4682 42464
rect 4618 42404 4622 42460
rect 4622 42404 4678 42460
rect 4678 42404 4682 42460
rect 4618 42400 4682 42404
rect 7805 42460 7869 42464
rect 7805 42404 7809 42460
rect 7809 42404 7865 42460
rect 7865 42404 7869 42460
rect 7805 42400 7869 42404
rect 7885 42460 7949 42464
rect 7885 42404 7889 42460
rect 7889 42404 7945 42460
rect 7945 42404 7949 42460
rect 7885 42400 7949 42404
rect 7965 42460 8029 42464
rect 7965 42404 7969 42460
rect 7969 42404 8025 42460
rect 8025 42404 8029 42460
rect 7965 42400 8029 42404
rect 8045 42460 8109 42464
rect 8045 42404 8049 42460
rect 8049 42404 8105 42460
rect 8105 42404 8109 42460
rect 8045 42400 8109 42404
rect 11232 42460 11296 42464
rect 11232 42404 11236 42460
rect 11236 42404 11292 42460
rect 11292 42404 11296 42460
rect 11232 42400 11296 42404
rect 11312 42460 11376 42464
rect 11312 42404 11316 42460
rect 11316 42404 11372 42460
rect 11372 42404 11376 42460
rect 11312 42400 11376 42404
rect 11392 42460 11456 42464
rect 11392 42404 11396 42460
rect 11396 42404 11452 42460
rect 11452 42404 11456 42460
rect 11392 42400 11456 42404
rect 11472 42460 11536 42464
rect 11472 42404 11476 42460
rect 11476 42404 11532 42460
rect 11532 42404 11536 42460
rect 11472 42400 11536 42404
rect 14659 42460 14723 42464
rect 14659 42404 14663 42460
rect 14663 42404 14719 42460
rect 14719 42404 14723 42460
rect 14659 42400 14723 42404
rect 14739 42460 14803 42464
rect 14739 42404 14743 42460
rect 14743 42404 14799 42460
rect 14799 42404 14803 42460
rect 14739 42400 14803 42404
rect 14819 42460 14883 42464
rect 14819 42404 14823 42460
rect 14823 42404 14879 42460
rect 14879 42404 14883 42460
rect 14819 42400 14883 42404
rect 14899 42460 14963 42464
rect 14899 42404 14903 42460
rect 14903 42404 14959 42460
rect 14959 42404 14963 42460
rect 14899 42400 14963 42404
rect 2665 41916 2729 41920
rect 2665 41860 2669 41916
rect 2669 41860 2725 41916
rect 2725 41860 2729 41916
rect 2665 41856 2729 41860
rect 2745 41916 2809 41920
rect 2745 41860 2749 41916
rect 2749 41860 2805 41916
rect 2805 41860 2809 41916
rect 2745 41856 2809 41860
rect 2825 41916 2889 41920
rect 2825 41860 2829 41916
rect 2829 41860 2885 41916
rect 2885 41860 2889 41916
rect 2825 41856 2889 41860
rect 2905 41916 2969 41920
rect 2905 41860 2909 41916
rect 2909 41860 2965 41916
rect 2965 41860 2969 41916
rect 2905 41856 2969 41860
rect 6092 41916 6156 41920
rect 6092 41860 6096 41916
rect 6096 41860 6152 41916
rect 6152 41860 6156 41916
rect 6092 41856 6156 41860
rect 6172 41916 6236 41920
rect 6172 41860 6176 41916
rect 6176 41860 6232 41916
rect 6232 41860 6236 41916
rect 6172 41856 6236 41860
rect 6252 41916 6316 41920
rect 6252 41860 6256 41916
rect 6256 41860 6312 41916
rect 6312 41860 6316 41916
rect 6252 41856 6316 41860
rect 6332 41916 6396 41920
rect 6332 41860 6336 41916
rect 6336 41860 6392 41916
rect 6392 41860 6396 41916
rect 6332 41856 6396 41860
rect 9519 41916 9583 41920
rect 9519 41860 9523 41916
rect 9523 41860 9579 41916
rect 9579 41860 9583 41916
rect 9519 41856 9583 41860
rect 9599 41916 9663 41920
rect 9599 41860 9603 41916
rect 9603 41860 9659 41916
rect 9659 41860 9663 41916
rect 9599 41856 9663 41860
rect 9679 41916 9743 41920
rect 9679 41860 9683 41916
rect 9683 41860 9739 41916
rect 9739 41860 9743 41916
rect 9679 41856 9743 41860
rect 9759 41916 9823 41920
rect 9759 41860 9763 41916
rect 9763 41860 9819 41916
rect 9819 41860 9823 41916
rect 9759 41856 9823 41860
rect 12946 41916 13010 41920
rect 12946 41860 12950 41916
rect 12950 41860 13006 41916
rect 13006 41860 13010 41916
rect 12946 41856 13010 41860
rect 13026 41916 13090 41920
rect 13026 41860 13030 41916
rect 13030 41860 13086 41916
rect 13086 41860 13090 41916
rect 13026 41856 13090 41860
rect 13106 41916 13170 41920
rect 13106 41860 13110 41916
rect 13110 41860 13166 41916
rect 13166 41860 13170 41916
rect 13106 41856 13170 41860
rect 13186 41916 13250 41920
rect 13186 41860 13190 41916
rect 13190 41860 13246 41916
rect 13246 41860 13250 41916
rect 13186 41856 13250 41860
rect 4378 41372 4442 41376
rect 4378 41316 4382 41372
rect 4382 41316 4438 41372
rect 4438 41316 4442 41372
rect 4378 41312 4442 41316
rect 4458 41372 4522 41376
rect 4458 41316 4462 41372
rect 4462 41316 4518 41372
rect 4518 41316 4522 41372
rect 4458 41312 4522 41316
rect 4538 41372 4602 41376
rect 4538 41316 4542 41372
rect 4542 41316 4598 41372
rect 4598 41316 4602 41372
rect 4538 41312 4602 41316
rect 4618 41372 4682 41376
rect 4618 41316 4622 41372
rect 4622 41316 4678 41372
rect 4678 41316 4682 41372
rect 4618 41312 4682 41316
rect 7805 41372 7869 41376
rect 7805 41316 7809 41372
rect 7809 41316 7865 41372
rect 7865 41316 7869 41372
rect 7805 41312 7869 41316
rect 7885 41372 7949 41376
rect 7885 41316 7889 41372
rect 7889 41316 7945 41372
rect 7945 41316 7949 41372
rect 7885 41312 7949 41316
rect 7965 41372 8029 41376
rect 7965 41316 7969 41372
rect 7969 41316 8025 41372
rect 8025 41316 8029 41372
rect 7965 41312 8029 41316
rect 8045 41372 8109 41376
rect 8045 41316 8049 41372
rect 8049 41316 8105 41372
rect 8105 41316 8109 41372
rect 8045 41312 8109 41316
rect 11232 41372 11296 41376
rect 11232 41316 11236 41372
rect 11236 41316 11292 41372
rect 11292 41316 11296 41372
rect 11232 41312 11296 41316
rect 11312 41372 11376 41376
rect 11312 41316 11316 41372
rect 11316 41316 11372 41372
rect 11372 41316 11376 41372
rect 11312 41312 11376 41316
rect 11392 41372 11456 41376
rect 11392 41316 11396 41372
rect 11396 41316 11452 41372
rect 11452 41316 11456 41372
rect 11392 41312 11456 41316
rect 11472 41372 11536 41376
rect 11472 41316 11476 41372
rect 11476 41316 11532 41372
rect 11532 41316 11536 41372
rect 11472 41312 11536 41316
rect 14659 41372 14723 41376
rect 14659 41316 14663 41372
rect 14663 41316 14719 41372
rect 14719 41316 14723 41372
rect 14659 41312 14723 41316
rect 14739 41372 14803 41376
rect 14739 41316 14743 41372
rect 14743 41316 14799 41372
rect 14799 41316 14803 41372
rect 14739 41312 14803 41316
rect 14819 41372 14883 41376
rect 14819 41316 14823 41372
rect 14823 41316 14879 41372
rect 14879 41316 14883 41372
rect 14819 41312 14883 41316
rect 14899 41372 14963 41376
rect 14899 41316 14903 41372
rect 14903 41316 14959 41372
rect 14959 41316 14963 41372
rect 14899 41312 14963 41316
rect 2665 40828 2729 40832
rect 2665 40772 2669 40828
rect 2669 40772 2725 40828
rect 2725 40772 2729 40828
rect 2665 40768 2729 40772
rect 2745 40828 2809 40832
rect 2745 40772 2749 40828
rect 2749 40772 2805 40828
rect 2805 40772 2809 40828
rect 2745 40768 2809 40772
rect 2825 40828 2889 40832
rect 2825 40772 2829 40828
rect 2829 40772 2885 40828
rect 2885 40772 2889 40828
rect 2825 40768 2889 40772
rect 2905 40828 2969 40832
rect 2905 40772 2909 40828
rect 2909 40772 2965 40828
rect 2965 40772 2969 40828
rect 2905 40768 2969 40772
rect 6092 40828 6156 40832
rect 6092 40772 6096 40828
rect 6096 40772 6152 40828
rect 6152 40772 6156 40828
rect 6092 40768 6156 40772
rect 6172 40828 6236 40832
rect 6172 40772 6176 40828
rect 6176 40772 6232 40828
rect 6232 40772 6236 40828
rect 6172 40768 6236 40772
rect 6252 40828 6316 40832
rect 6252 40772 6256 40828
rect 6256 40772 6312 40828
rect 6312 40772 6316 40828
rect 6252 40768 6316 40772
rect 6332 40828 6396 40832
rect 6332 40772 6336 40828
rect 6336 40772 6392 40828
rect 6392 40772 6396 40828
rect 6332 40768 6396 40772
rect 9519 40828 9583 40832
rect 9519 40772 9523 40828
rect 9523 40772 9579 40828
rect 9579 40772 9583 40828
rect 9519 40768 9583 40772
rect 9599 40828 9663 40832
rect 9599 40772 9603 40828
rect 9603 40772 9659 40828
rect 9659 40772 9663 40828
rect 9599 40768 9663 40772
rect 9679 40828 9743 40832
rect 9679 40772 9683 40828
rect 9683 40772 9739 40828
rect 9739 40772 9743 40828
rect 9679 40768 9743 40772
rect 9759 40828 9823 40832
rect 9759 40772 9763 40828
rect 9763 40772 9819 40828
rect 9819 40772 9823 40828
rect 9759 40768 9823 40772
rect 12946 40828 13010 40832
rect 12946 40772 12950 40828
rect 12950 40772 13006 40828
rect 13006 40772 13010 40828
rect 12946 40768 13010 40772
rect 13026 40828 13090 40832
rect 13026 40772 13030 40828
rect 13030 40772 13086 40828
rect 13086 40772 13090 40828
rect 13026 40768 13090 40772
rect 13106 40828 13170 40832
rect 13106 40772 13110 40828
rect 13110 40772 13166 40828
rect 13166 40772 13170 40828
rect 13106 40768 13170 40772
rect 13186 40828 13250 40832
rect 13186 40772 13190 40828
rect 13190 40772 13246 40828
rect 13246 40772 13250 40828
rect 13186 40768 13250 40772
rect 4378 40284 4442 40288
rect 4378 40228 4382 40284
rect 4382 40228 4438 40284
rect 4438 40228 4442 40284
rect 4378 40224 4442 40228
rect 4458 40284 4522 40288
rect 4458 40228 4462 40284
rect 4462 40228 4518 40284
rect 4518 40228 4522 40284
rect 4458 40224 4522 40228
rect 4538 40284 4602 40288
rect 4538 40228 4542 40284
rect 4542 40228 4598 40284
rect 4598 40228 4602 40284
rect 4538 40224 4602 40228
rect 4618 40284 4682 40288
rect 4618 40228 4622 40284
rect 4622 40228 4678 40284
rect 4678 40228 4682 40284
rect 4618 40224 4682 40228
rect 7805 40284 7869 40288
rect 7805 40228 7809 40284
rect 7809 40228 7865 40284
rect 7865 40228 7869 40284
rect 7805 40224 7869 40228
rect 7885 40284 7949 40288
rect 7885 40228 7889 40284
rect 7889 40228 7945 40284
rect 7945 40228 7949 40284
rect 7885 40224 7949 40228
rect 7965 40284 8029 40288
rect 7965 40228 7969 40284
rect 7969 40228 8025 40284
rect 8025 40228 8029 40284
rect 7965 40224 8029 40228
rect 8045 40284 8109 40288
rect 8045 40228 8049 40284
rect 8049 40228 8105 40284
rect 8105 40228 8109 40284
rect 8045 40224 8109 40228
rect 11232 40284 11296 40288
rect 11232 40228 11236 40284
rect 11236 40228 11292 40284
rect 11292 40228 11296 40284
rect 11232 40224 11296 40228
rect 11312 40284 11376 40288
rect 11312 40228 11316 40284
rect 11316 40228 11372 40284
rect 11372 40228 11376 40284
rect 11312 40224 11376 40228
rect 11392 40284 11456 40288
rect 11392 40228 11396 40284
rect 11396 40228 11452 40284
rect 11452 40228 11456 40284
rect 11392 40224 11456 40228
rect 11472 40284 11536 40288
rect 11472 40228 11476 40284
rect 11476 40228 11532 40284
rect 11532 40228 11536 40284
rect 11472 40224 11536 40228
rect 14659 40284 14723 40288
rect 14659 40228 14663 40284
rect 14663 40228 14719 40284
rect 14719 40228 14723 40284
rect 14659 40224 14723 40228
rect 14739 40284 14803 40288
rect 14739 40228 14743 40284
rect 14743 40228 14799 40284
rect 14799 40228 14803 40284
rect 14739 40224 14803 40228
rect 14819 40284 14883 40288
rect 14819 40228 14823 40284
rect 14823 40228 14879 40284
rect 14879 40228 14883 40284
rect 14819 40224 14883 40228
rect 14899 40284 14963 40288
rect 14899 40228 14903 40284
rect 14903 40228 14959 40284
rect 14959 40228 14963 40284
rect 14899 40224 14963 40228
rect 2665 39740 2729 39744
rect 2665 39684 2669 39740
rect 2669 39684 2725 39740
rect 2725 39684 2729 39740
rect 2665 39680 2729 39684
rect 2745 39740 2809 39744
rect 2745 39684 2749 39740
rect 2749 39684 2805 39740
rect 2805 39684 2809 39740
rect 2745 39680 2809 39684
rect 2825 39740 2889 39744
rect 2825 39684 2829 39740
rect 2829 39684 2885 39740
rect 2885 39684 2889 39740
rect 2825 39680 2889 39684
rect 2905 39740 2969 39744
rect 2905 39684 2909 39740
rect 2909 39684 2965 39740
rect 2965 39684 2969 39740
rect 2905 39680 2969 39684
rect 6092 39740 6156 39744
rect 6092 39684 6096 39740
rect 6096 39684 6152 39740
rect 6152 39684 6156 39740
rect 6092 39680 6156 39684
rect 6172 39740 6236 39744
rect 6172 39684 6176 39740
rect 6176 39684 6232 39740
rect 6232 39684 6236 39740
rect 6172 39680 6236 39684
rect 6252 39740 6316 39744
rect 6252 39684 6256 39740
rect 6256 39684 6312 39740
rect 6312 39684 6316 39740
rect 6252 39680 6316 39684
rect 6332 39740 6396 39744
rect 6332 39684 6336 39740
rect 6336 39684 6392 39740
rect 6392 39684 6396 39740
rect 6332 39680 6396 39684
rect 9519 39740 9583 39744
rect 9519 39684 9523 39740
rect 9523 39684 9579 39740
rect 9579 39684 9583 39740
rect 9519 39680 9583 39684
rect 9599 39740 9663 39744
rect 9599 39684 9603 39740
rect 9603 39684 9659 39740
rect 9659 39684 9663 39740
rect 9599 39680 9663 39684
rect 9679 39740 9743 39744
rect 9679 39684 9683 39740
rect 9683 39684 9739 39740
rect 9739 39684 9743 39740
rect 9679 39680 9743 39684
rect 9759 39740 9823 39744
rect 9759 39684 9763 39740
rect 9763 39684 9819 39740
rect 9819 39684 9823 39740
rect 9759 39680 9823 39684
rect 12946 39740 13010 39744
rect 12946 39684 12950 39740
rect 12950 39684 13006 39740
rect 13006 39684 13010 39740
rect 12946 39680 13010 39684
rect 13026 39740 13090 39744
rect 13026 39684 13030 39740
rect 13030 39684 13086 39740
rect 13086 39684 13090 39740
rect 13026 39680 13090 39684
rect 13106 39740 13170 39744
rect 13106 39684 13110 39740
rect 13110 39684 13166 39740
rect 13166 39684 13170 39740
rect 13106 39680 13170 39684
rect 13186 39740 13250 39744
rect 13186 39684 13190 39740
rect 13190 39684 13246 39740
rect 13246 39684 13250 39740
rect 13186 39680 13250 39684
rect 4378 39196 4442 39200
rect 4378 39140 4382 39196
rect 4382 39140 4438 39196
rect 4438 39140 4442 39196
rect 4378 39136 4442 39140
rect 4458 39196 4522 39200
rect 4458 39140 4462 39196
rect 4462 39140 4518 39196
rect 4518 39140 4522 39196
rect 4458 39136 4522 39140
rect 4538 39196 4602 39200
rect 4538 39140 4542 39196
rect 4542 39140 4598 39196
rect 4598 39140 4602 39196
rect 4538 39136 4602 39140
rect 4618 39196 4682 39200
rect 4618 39140 4622 39196
rect 4622 39140 4678 39196
rect 4678 39140 4682 39196
rect 4618 39136 4682 39140
rect 7805 39196 7869 39200
rect 7805 39140 7809 39196
rect 7809 39140 7865 39196
rect 7865 39140 7869 39196
rect 7805 39136 7869 39140
rect 7885 39196 7949 39200
rect 7885 39140 7889 39196
rect 7889 39140 7945 39196
rect 7945 39140 7949 39196
rect 7885 39136 7949 39140
rect 7965 39196 8029 39200
rect 7965 39140 7969 39196
rect 7969 39140 8025 39196
rect 8025 39140 8029 39196
rect 7965 39136 8029 39140
rect 8045 39196 8109 39200
rect 8045 39140 8049 39196
rect 8049 39140 8105 39196
rect 8105 39140 8109 39196
rect 8045 39136 8109 39140
rect 11232 39196 11296 39200
rect 11232 39140 11236 39196
rect 11236 39140 11292 39196
rect 11292 39140 11296 39196
rect 11232 39136 11296 39140
rect 11312 39196 11376 39200
rect 11312 39140 11316 39196
rect 11316 39140 11372 39196
rect 11372 39140 11376 39196
rect 11312 39136 11376 39140
rect 11392 39196 11456 39200
rect 11392 39140 11396 39196
rect 11396 39140 11452 39196
rect 11452 39140 11456 39196
rect 11392 39136 11456 39140
rect 11472 39196 11536 39200
rect 11472 39140 11476 39196
rect 11476 39140 11532 39196
rect 11532 39140 11536 39196
rect 11472 39136 11536 39140
rect 14659 39196 14723 39200
rect 14659 39140 14663 39196
rect 14663 39140 14719 39196
rect 14719 39140 14723 39196
rect 14659 39136 14723 39140
rect 14739 39196 14803 39200
rect 14739 39140 14743 39196
rect 14743 39140 14799 39196
rect 14799 39140 14803 39196
rect 14739 39136 14803 39140
rect 14819 39196 14883 39200
rect 14819 39140 14823 39196
rect 14823 39140 14879 39196
rect 14879 39140 14883 39196
rect 14819 39136 14883 39140
rect 14899 39196 14963 39200
rect 14899 39140 14903 39196
rect 14903 39140 14959 39196
rect 14959 39140 14963 39196
rect 14899 39136 14963 39140
rect 2665 38652 2729 38656
rect 2665 38596 2669 38652
rect 2669 38596 2725 38652
rect 2725 38596 2729 38652
rect 2665 38592 2729 38596
rect 2745 38652 2809 38656
rect 2745 38596 2749 38652
rect 2749 38596 2805 38652
rect 2805 38596 2809 38652
rect 2745 38592 2809 38596
rect 2825 38652 2889 38656
rect 2825 38596 2829 38652
rect 2829 38596 2885 38652
rect 2885 38596 2889 38652
rect 2825 38592 2889 38596
rect 2905 38652 2969 38656
rect 2905 38596 2909 38652
rect 2909 38596 2965 38652
rect 2965 38596 2969 38652
rect 2905 38592 2969 38596
rect 6092 38652 6156 38656
rect 6092 38596 6096 38652
rect 6096 38596 6152 38652
rect 6152 38596 6156 38652
rect 6092 38592 6156 38596
rect 6172 38652 6236 38656
rect 6172 38596 6176 38652
rect 6176 38596 6232 38652
rect 6232 38596 6236 38652
rect 6172 38592 6236 38596
rect 6252 38652 6316 38656
rect 6252 38596 6256 38652
rect 6256 38596 6312 38652
rect 6312 38596 6316 38652
rect 6252 38592 6316 38596
rect 6332 38652 6396 38656
rect 6332 38596 6336 38652
rect 6336 38596 6392 38652
rect 6392 38596 6396 38652
rect 6332 38592 6396 38596
rect 9519 38652 9583 38656
rect 9519 38596 9523 38652
rect 9523 38596 9579 38652
rect 9579 38596 9583 38652
rect 9519 38592 9583 38596
rect 9599 38652 9663 38656
rect 9599 38596 9603 38652
rect 9603 38596 9659 38652
rect 9659 38596 9663 38652
rect 9599 38592 9663 38596
rect 9679 38652 9743 38656
rect 9679 38596 9683 38652
rect 9683 38596 9739 38652
rect 9739 38596 9743 38652
rect 9679 38592 9743 38596
rect 9759 38652 9823 38656
rect 9759 38596 9763 38652
rect 9763 38596 9819 38652
rect 9819 38596 9823 38652
rect 9759 38592 9823 38596
rect 12946 38652 13010 38656
rect 12946 38596 12950 38652
rect 12950 38596 13006 38652
rect 13006 38596 13010 38652
rect 12946 38592 13010 38596
rect 13026 38652 13090 38656
rect 13026 38596 13030 38652
rect 13030 38596 13086 38652
rect 13086 38596 13090 38652
rect 13026 38592 13090 38596
rect 13106 38652 13170 38656
rect 13106 38596 13110 38652
rect 13110 38596 13166 38652
rect 13166 38596 13170 38652
rect 13106 38592 13170 38596
rect 13186 38652 13250 38656
rect 13186 38596 13190 38652
rect 13190 38596 13246 38652
rect 13246 38596 13250 38652
rect 13186 38592 13250 38596
rect 4378 38108 4442 38112
rect 4378 38052 4382 38108
rect 4382 38052 4438 38108
rect 4438 38052 4442 38108
rect 4378 38048 4442 38052
rect 4458 38108 4522 38112
rect 4458 38052 4462 38108
rect 4462 38052 4518 38108
rect 4518 38052 4522 38108
rect 4458 38048 4522 38052
rect 4538 38108 4602 38112
rect 4538 38052 4542 38108
rect 4542 38052 4598 38108
rect 4598 38052 4602 38108
rect 4538 38048 4602 38052
rect 4618 38108 4682 38112
rect 4618 38052 4622 38108
rect 4622 38052 4678 38108
rect 4678 38052 4682 38108
rect 4618 38048 4682 38052
rect 7805 38108 7869 38112
rect 7805 38052 7809 38108
rect 7809 38052 7865 38108
rect 7865 38052 7869 38108
rect 7805 38048 7869 38052
rect 7885 38108 7949 38112
rect 7885 38052 7889 38108
rect 7889 38052 7945 38108
rect 7945 38052 7949 38108
rect 7885 38048 7949 38052
rect 7965 38108 8029 38112
rect 7965 38052 7969 38108
rect 7969 38052 8025 38108
rect 8025 38052 8029 38108
rect 7965 38048 8029 38052
rect 8045 38108 8109 38112
rect 8045 38052 8049 38108
rect 8049 38052 8105 38108
rect 8105 38052 8109 38108
rect 8045 38048 8109 38052
rect 11232 38108 11296 38112
rect 11232 38052 11236 38108
rect 11236 38052 11292 38108
rect 11292 38052 11296 38108
rect 11232 38048 11296 38052
rect 11312 38108 11376 38112
rect 11312 38052 11316 38108
rect 11316 38052 11372 38108
rect 11372 38052 11376 38108
rect 11312 38048 11376 38052
rect 11392 38108 11456 38112
rect 11392 38052 11396 38108
rect 11396 38052 11452 38108
rect 11452 38052 11456 38108
rect 11392 38048 11456 38052
rect 11472 38108 11536 38112
rect 11472 38052 11476 38108
rect 11476 38052 11532 38108
rect 11532 38052 11536 38108
rect 11472 38048 11536 38052
rect 14659 38108 14723 38112
rect 14659 38052 14663 38108
rect 14663 38052 14719 38108
rect 14719 38052 14723 38108
rect 14659 38048 14723 38052
rect 14739 38108 14803 38112
rect 14739 38052 14743 38108
rect 14743 38052 14799 38108
rect 14799 38052 14803 38108
rect 14739 38048 14803 38052
rect 14819 38108 14883 38112
rect 14819 38052 14823 38108
rect 14823 38052 14879 38108
rect 14879 38052 14883 38108
rect 14819 38048 14883 38052
rect 14899 38108 14963 38112
rect 14899 38052 14903 38108
rect 14903 38052 14959 38108
rect 14959 38052 14963 38108
rect 14899 38048 14963 38052
rect 2665 37564 2729 37568
rect 2665 37508 2669 37564
rect 2669 37508 2725 37564
rect 2725 37508 2729 37564
rect 2665 37504 2729 37508
rect 2745 37564 2809 37568
rect 2745 37508 2749 37564
rect 2749 37508 2805 37564
rect 2805 37508 2809 37564
rect 2745 37504 2809 37508
rect 2825 37564 2889 37568
rect 2825 37508 2829 37564
rect 2829 37508 2885 37564
rect 2885 37508 2889 37564
rect 2825 37504 2889 37508
rect 2905 37564 2969 37568
rect 2905 37508 2909 37564
rect 2909 37508 2965 37564
rect 2965 37508 2969 37564
rect 2905 37504 2969 37508
rect 6092 37564 6156 37568
rect 6092 37508 6096 37564
rect 6096 37508 6152 37564
rect 6152 37508 6156 37564
rect 6092 37504 6156 37508
rect 6172 37564 6236 37568
rect 6172 37508 6176 37564
rect 6176 37508 6232 37564
rect 6232 37508 6236 37564
rect 6172 37504 6236 37508
rect 6252 37564 6316 37568
rect 6252 37508 6256 37564
rect 6256 37508 6312 37564
rect 6312 37508 6316 37564
rect 6252 37504 6316 37508
rect 6332 37564 6396 37568
rect 6332 37508 6336 37564
rect 6336 37508 6392 37564
rect 6392 37508 6396 37564
rect 6332 37504 6396 37508
rect 9519 37564 9583 37568
rect 9519 37508 9523 37564
rect 9523 37508 9579 37564
rect 9579 37508 9583 37564
rect 9519 37504 9583 37508
rect 9599 37564 9663 37568
rect 9599 37508 9603 37564
rect 9603 37508 9659 37564
rect 9659 37508 9663 37564
rect 9599 37504 9663 37508
rect 9679 37564 9743 37568
rect 9679 37508 9683 37564
rect 9683 37508 9739 37564
rect 9739 37508 9743 37564
rect 9679 37504 9743 37508
rect 9759 37564 9823 37568
rect 9759 37508 9763 37564
rect 9763 37508 9819 37564
rect 9819 37508 9823 37564
rect 9759 37504 9823 37508
rect 12946 37564 13010 37568
rect 12946 37508 12950 37564
rect 12950 37508 13006 37564
rect 13006 37508 13010 37564
rect 12946 37504 13010 37508
rect 13026 37564 13090 37568
rect 13026 37508 13030 37564
rect 13030 37508 13086 37564
rect 13086 37508 13090 37564
rect 13026 37504 13090 37508
rect 13106 37564 13170 37568
rect 13106 37508 13110 37564
rect 13110 37508 13166 37564
rect 13166 37508 13170 37564
rect 13106 37504 13170 37508
rect 13186 37564 13250 37568
rect 13186 37508 13190 37564
rect 13190 37508 13246 37564
rect 13246 37508 13250 37564
rect 13186 37504 13250 37508
rect 4378 37020 4442 37024
rect 4378 36964 4382 37020
rect 4382 36964 4438 37020
rect 4438 36964 4442 37020
rect 4378 36960 4442 36964
rect 4458 37020 4522 37024
rect 4458 36964 4462 37020
rect 4462 36964 4518 37020
rect 4518 36964 4522 37020
rect 4458 36960 4522 36964
rect 4538 37020 4602 37024
rect 4538 36964 4542 37020
rect 4542 36964 4598 37020
rect 4598 36964 4602 37020
rect 4538 36960 4602 36964
rect 4618 37020 4682 37024
rect 4618 36964 4622 37020
rect 4622 36964 4678 37020
rect 4678 36964 4682 37020
rect 4618 36960 4682 36964
rect 7805 37020 7869 37024
rect 7805 36964 7809 37020
rect 7809 36964 7865 37020
rect 7865 36964 7869 37020
rect 7805 36960 7869 36964
rect 7885 37020 7949 37024
rect 7885 36964 7889 37020
rect 7889 36964 7945 37020
rect 7945 36964 7949 37020
rect 7885 36960 7949 36964
rect 7965 37020 8029 37024
rect 7965 36964 7969 37020
rect 7969 36964 8025 37020
rect 8025 36964 8029 37020
rect 7965 36960 8029 36964
rect 8045 37020 8109 37024
rect 8045 36964 8049 37020
rect 8049 36964 8105 37020
rect 8105 36964 8109 37020
rect 8045 36960 8109 36964
rect 11232 37020 11296 37024
rect 11232 36964 11236 37020
rect 11236 36964 11292 37020
rect 11292 36964 11296 37020
rect 11232 36960 11296 36964
rect 11312 37020 11376 37024
rect 11312 36964 11316 37020
rect 11316 36964 11372 37020
rect 11372 36964 11376 37020
rect 11312 36960 11376 36964
rect 11392 37020 11456 37024
rect 11392 36964 11396 37020
rect 11396 36964 11452 37020
rect 11452 36964 11456 37020
rect 11392 36960 11456 36964
rect 11472 37020 11536 37024
rect 11472 36964 11476 37020
rect 11476 36964 11532 37020
rect 11532 36964 11536 37020
rect 11472 36960 11536 36964
rect 14659 37020 14723 37024
rect 14659 36964 14663 37020
rect 14663 36964 14719 37020
rect 14719 36964 14723 37020
rect 14659 36960 14723 36964
rect 14739 37020 14803 37024
rect 14739 36964 14743 37020
rect 14743 36964 14799 37020
rect 14799 36964 14803 37020
rect 14739 36960 14803 36964
rect 14819 37020 14883 37024
rect 14819 36964 14823 37020
rect 14823 36964 14879 37020
rect 14879 36964 14883 37020
rect 14819 36960 14883 36964
rect 14899 37020 14963 37024
rect 14899 36964 14903 37020
rect 14903 36964 14959 37020
rect 14959 36964 14963 37020
rect 14899 36960 14963 36964
rect 2665 36476 2729 36480
rect 2665 36420 2669 36476
rect 2669 36420 2725 36476
rect 2725 36420 2729 36476
rect 2665 36416 2729 36420
rect 2745 36476 2809 36480
rect 2745 36420 2749 36476
rect 2749 36420 2805 36476
rect 2805 36420 2809 36476
rect 2745 36416 2809 36420
rect 2825 36476 2889 36480
rect 2825 36420 2829 36476
rect 2829 36420 2885 36476
rect 2885 36420 2889 36476
rect 2825 36416 2889 36420
rect 2905 36476 2969 36480
rect 2905 36420 2909 36476
rect 2909 36420 2965 36476
rect 2965 36420 2969 36476
rect 2905 36416 2969 36420
rect 6092 36476 6156 36480
rect 6092 36420 6096 36476
rect 6096 36420 6152 36476
rect 6152 36420 6156 36476
rect 6092 36416 6156 36420
rect 6172 36476 6236 36480
rect 6172 36420 6176 36476
rect 6176 36420 6232 36476
rect 6232 36420 6236 36476
rect 6172 36416 6236 36420
rect 6252 36476 6316 36480
rect 6252 36420 6256 36476
rect 6256 36420 6312 36476
rect 6312 36420 6316 36476
rect 6252 36416 6316 36420
rect 6332 36476 6396 36480
rect 6332 36420 6336 36476
rect 6336 36420 6392 36476
rect 6392 36420 6396 36476
rect 6332 36416 6396 36420
rect 9519 36476 9583 36480
rect 9519 36420 9523 36476
rect 9523 36420 9579 36476
rect 9579 36420 9583 36476
rect 9519 36416 9583 36420
rect 9599 36476 9663 36480
rect 9599 36420 9603 36476
rect 9603 36420 9659 36476
rect 9659 36420 9663 36476
rect 9599 36416 9663 36420
rect 9679 36476 9743 36480
rect 9679 36420 9683 36476
rect 9683 36420 9739 36476
rect 9739 36420 9743 36476
rect 9679 36416 9743 36420
rect 9759 36476 9823 36480
rect 9759 36420 9763 36476
rect 9763 36420 9819 36476
rect 9819 36420 9823 36476
rect 9759 36416 9823 36420
rect 12946 36476 13010 36480
rect 12946 36420 12950 36476
rect 12950 36420 13006 36476
rect 13006 36420 13010 36476
rect 12946 36416 13010 36420
rect 13026 36476 13090 36480
rect 13026 36420 13030 36476
rect 13030 36420 13086 36476
rect 13086 36420 13090 36476
rect 13026 36416 13090 36420
rect 13106 36476 13170 36480
rect 13106 36420 13110 36476
rect 13110 36420 13166 36476
rect 13166 36420 13170 36476
rect 13106 36416 13170 36420
rect 13186 36476 13250 36480
rect 13186 36420 13190 36476
rect 13190 36420 13246 36476
rect 13246 36420 13250 36476
rect 13186 36416 13250 36420
rect 4378 35932 4442 35936
rect 4378 35876 4382 35932
rect 4382 35876 4438 35932
rect 4438 35876 4442 35932
rect 4378 35872 4442 35876
rect 4458 35932 4522 35936
rect 4458 35876 4462 35932
rect 4462 35876 4518 35932
rect 4518 35876 4522 35932
rect 4458 35872 4522 35876
rect 4538 35932 4602 35936
rect 4538 35876 4542 35932
rect 4542 35876 4598 35932
rect 4598 35876 4602 35932
rect 4538 35872 4602 35876
rect 4618 35932 4682 35936
rect 4618 35876 4622 35932
rect 4622 35876 4678 35932
rect 4678 35876 4682 35932
rect 4618 35872 4682 35876
rect 7805 35932 7869 35936
rect 7805 35876 7809 35932
rect 7809 35876 7865 35932
rect 7865 35876 7869 35932
rect 7805 35872 7869 35876
rect 7885 35932 7949 35936
rect 7885 35876 7889 35932
rect 7889 35876 7945 35932
rect 7945 35876 7949 35932
rect 7885 35872 7949 35876
rect 7965 35932 8029 35936
rect 7965 35876 7969 35932
rect 7969 35876 8025 35932
rect 8025 35876 8029 35932
rect 7965 35872 8029 35876
rect 8045 35932 8109 35936
rect 8045 35876 8049 35932
rect 8049 35876 8105 35932
rect 8105 35876 8109 35932
rect 8045 35872 8109 35876
rect 11232 35932 11296 35936
rect 11232 35876 11236 35932
rect 11236 35876 11292 35932
rect 11292 35876 11296 35932
rect 11232 35872 11296 35876
rect 11312 35932 11376 35936
rect 11312 35876 11316 35932
rect 11316 35876 11372 35932
rect 11372 35876 11376 35932
rect 11312 35872 11376 35876
rect 11392 35932 11456 35936
rect 11392 35876 11396 35932
rect 11396 35876 11452 35932
rect 11452 35876 11456 35932
rect 11392 35872 11456 35876
rect 11472 35932 11536 35936
rect 11472 35876 11476 35932
rect 11476 35876 11532 35932
rect 11532 35876 11536 35932
rect 11472 35872 11536 35876
rect 14659 35932 14723 35936
rect 14659 35876 14663 35932
rect 14663 35876 14719 35932
rect 14719 35876 14723 35932
rect 14659 35872 14723 35876
rect 14739 35932 14803 35936
rect 14739 35876 14743 35932
rect 14743 35876 14799 35932
rect 14799 35876 14803 35932
rect 14739 35872 14803 35876
rect 14819 35932 14883 35936
rect 14819 35876 14823 35932
rect 14823 35876 14879 35932
rect 14879 35876 14883 35932
rect 14819 35872 14883 35876
rect 14899 35932 14963 35936
rect 14899 35876 14903 35932
rect 14903 35876 14959 35932
rect 14959 35876 14963 35932
rect 14899 35872 14963 35876
rect 2665 35388 2729 35392
rect 2665 35332 2669 35388
rect 2669 35332 2725 35388
rect 2725 35332 2729 35388
rect 2665 35328 2729 35332
rect 2745 35388 2809 35392
rect 2745 35332 2749 35388
rect 2749 35332 2805 35388
rect 2805 35332 2809 35388
rect 2745 35328 2809 35332
rect 2825 35388 2889 35392
rect 2825 35332 2829 35388
rect 2829 35332 2885 35388
rect 2885 35332 2889 35388
rect 2825 35328 2889 35332
rect 2905 35388 2969 35392
rect 2905 35332 2909 35388
rect 2909 35332 2965 35388
rect 2965 35332 2969 35388
rect 2905 35328 2969 35332
rect 6092 35388 6156 35392
rect 6092 35332 6096 35388
rect 6096 35332 6152 35388
rect 6152 35332 6156 35388
rect 6092 35328 6156 35332
rect 6172 35388 6236 35392
rect 6172 35332 6176 35388
rect 6176 35332 6232 35388
rect 6232 35332 6236 35388
rect 6172 35328 6236 35332
rect 6252 35388 6316 35392
rect 6252 35332 6256 35388
rect 6256 35332 6312 35388
rect 6312 35332 6316 35388
rect 6252 35328 6316 35332
rect 6332 35388 6396 35392
rect 6332 35332 6336 35388
rect 6336 35332 6392 35388
rect 6392 35332 6396 35388
rect 6332 35328 6396 35332
rect 9519 35388 9583 35392
rect 9519 35332 9523 35388
rect 9523 35332 9579 35388
rect 9579 35332 9583 35388
rect 9519 35328 9583 35332
rect 9599 35388 9663 35392
rect 9599 35332 9603 35388
rect 9603 35332 9659 35388
rect 9659 35332 9663 35388
rect 9599 35328 9663 35332
rect 9679 35388 9743 35392
rect 9679 35332 9683 35388
rect 9683 35332 9739 35388
rect 9739 35332 9743 35388
rect 9679 35328 9743 35332
rect 9759 35388 9823 35392
rect 9759 35332 9763 35388
rect 9763 35332 9819 35388
rect 9819 35332 9823 35388
rect 9759 35328 9823 35332
rect 12946 35388 13010 35392
rect 12946 35332 12950 35388
rect 12950 35332 13006 35388
rect 13006 35332 13010 35388
rect 12946 35328 13010 35332
rect 13026 35388 13090 35392
rect 13026 35332 13030 35388
rect 13030 35332 13086 35388
rect 13086 35332 13090 35388
rect 13026 35328 13090 35332
rect 13106 35388 13170 35392
rect 13106 35332 13110 35388
rect 13110 35332 13166 35388
rect 13166 35332 13170 35388
rect 13106 35328 13170 35332
rect 13186 35388 13250 35392
rect 13186 35332 13190 35388
rect 13190 35332 13246 35388
rect 13246 35332 13250 35388
rect 13186 35328 13250 35332
rect 4378 34844 4442 34848
rect 4378 34788 4382 34844
rect 4382 34788 4438 34844
rect 4438 34788 4442 34844
rect 4378 34784 4442 34788
rect 4458 34844 4522 34848
rect 4458 34788 4462 34844
rect 4462 34788 4518 34844
rect 4518 34788 4522 34844
rect 4458 34784 4522 34788
rect 4538 34844 4602 34848
rect 4538 34788 4542 34844
rect 4542 34788 4598 34844
rect 4598 34788 4602 34844
rect 4538 34784 4602 34788
rect 4618 34844 4682 34848
rect 4618 34788 4622 34844
rect 4622 34788 4678 34844
rect 4678 34788 4682 34844
rect 4618 34784 4682 34788
rect 7805 34844 7869 34848
rect 7805 34788 7809 34844
rect 7809 34788 7865 34844
rect 7865 34788 7869 34844
rect 7805 34784 7869 34788
rect 7885 34844 7949 34848
rect 7885 34788 7889 34844
rect 7889 34788 7945 34844
rect 7945 34788 7949 34844
rect 7885 34784 7949 34788
rect 7965 34844 8029 34848
rect 7965 34788 7969 34844
rect 7969 34788 8025 34844
rect 8025 34788 8029 34844
rect 7965 34784 8029 34788
rect 8045 34844 8109 34848
rect 8045 34788 8049 34844
rect 8049 34788 8105 34844
rect 8105 34788 8109 34844
rect 8045 34784 8109 34788
rect 11232 34844 11296 34848
rect 11232 34788 11236 34844
rect 11236 34788 11292 34844
rect 11292 34788 11296 34844
rect 11232 34784 11296 34788
rect 11312 34844 11376 34848
rect 11312 34788 11316 34844
rect 11316 34788 11372 34844
rect 11372 34788 11376 34844
rect 11312 34784 11376 34788
rect 11392 34844 11456 34848
rect 11392 34788 11396 34844
rect 11396 34788 11452 34844
rect 11452 34788 11456 34844
rect 11392 34784 11456 34788
rect 11472 34844 11536 34848
rect 11472 34788 11476 34844
rect 11476 34788 11532 34844
rect 11532 34788 11536 34844
rect 11472 34784 11536 34788
rect 14659 34844 14723 34848
rect 14659 34788 14663 34844
rect 14663 34788 14719 34844
rect 14719 34788 14723 34844
rect 14659 34784 14723 34788
rect 14739 34844 14803 34848
rect 14739 34788 14743 34844
rect 14743 34788 14799 34844
rect 14799 34788 14803 34844
rect 14739 34784 14803 34788
rect 14819 34844 14883 34848
rect 14819 34788 14823 34844
rect 14823 34788 14879 34844
rect 14879 34788 14883 34844
rect 14819 34784 14883 34788
rect 14899 34844 14963 34848
rect 14899 34788 14903 34844
rect 14903 34788 14959 34844
rect 14959 34788 14963 34844
rect 14899 34784 14963 34788
rect 2665 34300 2729 34304
rect 2665 34244 2669 34300
rect 2669 34244 2725 34300
rect 2725 34244 2729 34300
rect 2665 34240 2729 34244
rect 2745 34300 2809 34304
rect 2745 34244 2749 34300
rect 2749 34244 2805 34300
rect 2805 34244 2809 34300
rect 2745 34240 2809 34244
rect 2825 34300 2889 34304
rect 2825 34244 2829 34300
rect 2829 34244 2885 34300
rect 2885 34244 2889 34300
rect 2825 34240 2889 34244
rect 2905 34300 2969 34304
rect 2905 34244 2909 34300
rect 2909 34244 2965 34300
rect 2965 34244 2969 34300
rect 2905 34240 2969 34244
rect 6092 34300 6156 34304
rect 6092 34244 6096 34300
rect 6096 34244 6152 34300
rect 6152 34244 6156 34300
rect 6092 34240 6156 34244
rect 6172 34300 6236 34304
rect 6172 34244 6176 34300
rect 6176 34244 6232 34300
rect 6232 34244 6236 34300
rect 6172 34240 6236 34244
rect 6252 34300 6316 34304
rect 6252 34244 6256 34300
rect 6256 34244 6312 34300
rect 6312 34244 6316 34300
rect 6252 34240 6316 34244
rect 6332 34300 6396 34304
rect 6332 34244 6336 34300
rect 6336 34244 6392 34300
rect 6392 34244 6396 34300
rect 6332 34240 6396 34244
rect 9519 34300 9583 34304
rect 9519 34244 9523 34300
rect 9523 34244 9579 34300
rect 9579 34244 9583 34300
rect 9519 34240 9583 34244
rect 9599 34300 9663 34304
rect 9599 34244 9603 34300
rect 9603 34244 9659 34300
rect 9659 34244 9663 34300
rect 9599 34240 9663 34244
rect 9679 34300 9743 34304
rect 9679 34244 9683 34300
rect 9683 34244 9739 34300
rect 9739 34244 9743 34300
rect 9679 34240 9743 34244
rect 9759 34300 9823 34304
rect 9759 34244 9763 34300
rect 9763 34244 9819 34300
rect 9819 34244 9823 34300
rect 9759 34240 9823 34244
rect 12946 34300 13010 34304
rect 12946 34244 12950 34300
rect 12950 34244 13006 34300
rect 13006 34244 13010 34300
rect 12946 34240 13010 34244
rect 13026 34300 13090 34304
rect 13026 34244 13030 34300
rect 13030 34244 13086 34300
rect 13086 34244 13090 34300
rect 13026 34240 13090 34244
rect 13106 34300 13170 34304
rect 13106 34244 13110 34300
rect 13110 34244 13166 34300
rect 13166 34244 13170 34300
rect 13106 34240 13170 34244
rect 13186 34300 13250 34304
rect 13186 34244 13190 34300
rect 13190 34244 13246 34300
rect 13246 34244 13250 34300
rect 13186 34240 13250 34244
rect 4378 33756 4442 33760
rect 4378 33700 4382 33756
rect 4382 33700 4438 33756
rect 4438 33700 4442 33756
rect 4378 33696 4442 33700
rect 4458 33756 4522 33760
rect 4458 33700 4462 33756
rect 4462 33700 4518 33756
rect 4518 33700 4522 33756
rect 4458 33696 4522 33700
rect 4538 33756 4602 33760
rect 4538 33700 4542 33756
rect 4542 33700 4598 33756
rect 4598 33700 4602 33756
rect 4538 33696 4602 33700
rect 4618 33756 4682 33760
rect 4618 33700 4622 33756
rect 4622 33700 4678 33756
rect 4678 33700 4682 33756
rect 4618 33696 4682 33700
rect 7805 33756 7869 33760
rect 7805 33700 7809 33756
rect 7809 33700 7865 33756
rect 7865 33700 7869 33756
rect 7805 33696 7869 33700
rect 7885 33756 7949 33760
rect 7885 33700 7889 33756
rect 7889 33700 7945 33756
rect 7945 33700 7949 33756
rect 7885 33696 7949 33700
rect 7965 33756 8029 33760
rect 7965 33700 7969 33756
rect 7969 33700 8025 33756
rect 8025 33700 8029 33756
rect 7965 33696 8029 33700
rect 8045 33756 8109 33760
rect 8045 33700 8049 33756
rect 8049 33700 8105 33756
rect 8105 33700 8109 33756
rect 8045 33696 8109 33700
rect 11232 33756 11296 33760
rect 11232 33700 11236 33756
rect 11236 33700 11292 33756
rect 11292 33700 11296 33756
rect 11232 33696 11296 33700
rect 11312 33756 11376 33760
rect 11312 33700 11316 33756
rect 11316 33700 11372 33756
rect 11372 33700 11376 33756
rect 11312 33696 11376 33700
rect 11392 33756 11456 33760
rect 11392 33700 11396 33756
rect 11396 33700 11452 33756
rect 11452 33700 11456 33756
rect 11392 33696 11456 33700
rect 11472 33756 11536 33760
rect 11472 33700 11476 33756
rect 11476 33700 11532 33756
rect 11532 33700 11536 33756
rect 11472 33696 11536 33700
rect 14659 33756 14723 33760
rect 14659 33700 14663 33756
rect 14663 33700 14719 33756
rect 14719 33700 14723 33756
rect 14659 33696 14723 33700
rect 14739 33756 14803 33760
rect 14739 33700 14743 33756
rect 14743 33700 14799 33756
rect 14799 33700 14803 33756
rect 14739 33696 14803 33700
rect 14819 33756 14883 33760
rect 14819 33700 14823 33756
rect 14823 33700 14879 33756
rect 14879 33700 14883 33756
rect 14819 33696 14883 33700
rect 14899 33756 14963 33760
rect 14899 33700 14903 33756
rect 14903 33700 14959 33756
rect 14959 33700 14963 33756
rect 14899 33696 14963 33700
rect 2665 33212 2729 33216
rect 2665 33156 2669 33212
rect 2669 33156 2725 33212
rect 2725 33156 2729 33212
rect 2665 33152 2729 33156
rect 2745 33212 2809 33216
rect 2745 33156 2749 33212
rect 2749 33156 2805 33212
rect 2805 33156 2809 33212
rect 2745 33152 2809 33156
rect 2825 33212 2889 33216
rect 2825 33156 2829 33212
rect 2829 33156 2885 33212
rect 2885 33156 2889 33212
rect 2825 33152 2889 33156
rect 2905 33212 2969 33216
rect 2905 33156 2909 33212
rect 2909 33156 2965 33212
rect 2965 33156 2969 33212
rect 2905 33152 2969 33156
rect 6092 33212 6156 33216
rect 6092 33156 6096 33212
rect 6096 33156 6152 33212
rect 6152 33156 6156 33212
rect 6092 33152 6156 33156
rect 6172 33212 6236 33216
rect 6172 33156 6176 33212
rect 6176 33156 6232 33212
rect 6232 33156 6236 33212
rect 6172 33152 6236 33156
rect 6252 33212 6316 33216
rect 6252 33156 6256 33212
rect 6256 33156 6312 33212
rect 6312 33156 6316 33212
rect 6252 33152 6316 33156
rect 6332 33212 6396 33216
rect 6332 33156 6336 33212
rect 6336 33156 6392 33212
rect 6392 33156 6396 33212
rect 6332 33152 6396 33156
rect 9519 33212 9583 33216
rect 9519 33156 9523 33212
rect 9523 33156 9579 33212
rect 9579 33156 9583 33212
rect 9519 33152 9583 33156
rect 9599 33212 9663 33216
rect 9599 33156 9603 33212
rect 9603 33156 9659 33212
rect 9659 33156 9663 33212
rect 9599 33152 9663 33156
rect 9679 33212 9743 33216
rect 9679 33156 9683 33212
rect 9683 33156 9739 33212
rect 9739 33156 9743 33212
rect 9679 33152 9743 33156
rect 9759 33212 9823 33216
rect 9759 33156 9763 33212
rect 9763 33156 9819 33212
rect 9819 33156 9823 33212
rect 9759 33152 9823 33156
rect 12946 33212 13010 33216
rect 12946 33156 12950 33212
rect 12950 33156 13006 33212
rect 13006 33156 13010 33212
rect 12946 33152 13010 33156
rect 13026 33212 13090 33216
rect 13026 33156 13030 33212
rect 13030 33156 13086 33212
rect 13086 33156 13090 33212
rect 13026 33152 13090 33156
rect 13106 33212 13170 33216
rect 13106 33156 13110 33212
rect 13110 33156 13166 33212
rect 13166 33156 13170 33212
rect 13106 33152 13170 33156
rect 13186 33212 13250 33216
rect 13186 33156 13190 33212
rect 13190 33156 13246 33212
rect 13246 33156 13250 33212
rect 13186 33152 13250 33156
rect 4378 32668 4442 32672
rect 4378 32612 4382 32668
rect 4382 32612 4438 32668
rect 4438 32612 4442 32668
rect 4378 32608 4442 32612
rect 4458 32668 4522 32672
rect 4458 32612 4462 32668
rect 4462 32612 4518 32668
rect 4518 32612 4522 32668
rect 4458 32608 4522 32612
rect 4538 32668 4602 32672
rect 4538 32612 4542 32668
rect 4542 32612 4598 32668
rect 4598 32612 4602 32668
rect 4538 32608 4602 32612
rect 4618 32668 4682 32672
rect 4618 32612 4622 32668
rect 4622 32612 4678 32668
rect 4678 32612 4682 32668
rect 4618 32608 4682 32612
rect 7805 32668 7869 32672
rect 7805 32612 7809 32668
rect 7809 32612 7865 32668
rect 7865 32612 7869 32668
rect 7805 32608 7869 32612
rect 7885 32668 7949 32672
rect 7885 32612 7889 32668
rect 7889 32612 7945 32668
rect 7945 32612 7949 32668
rect 7885 32608 7949 32612
rect 7965 32668 8029 32672
rect 7965 32612 7969 32668
rect 7969 32612 8025 32668
rect 8025 32612 8029 32668
rect 7965 32608 8029 32612
rect 8045 32668 8109 32672
rect 8045 32612 8049 32668
rect 8049 32612 8105 32668
rect 8105 32612 8109 32668
rect 8045 32608 8109 32612
rect 11232 32668 11296 32672
rect 11232 32612 11236 32668
rect 11236 32612 11292 32668
rect 11292 32612 11296 32668
rect 11232 32608 11296 32612
rect 11312 32668 11376 32672
rect 11312 32612 11316 32668
rect 11316 32612 11372 32668
rect 11372 32612 11376 32668
rect 11312 32608 11376 32612
rect 11392 32668 11456 32672
rect 11392 32612 11396 32668
rect 11396 32612 11452 32668
rect 11452 32612 11456 32668
rect 11392 32608 11456 32612
rect 11472 32668 11536 32672
rect 11472 32612 11476 32668
rect 11476 32612 11532 32668
rect 11532 32612 11536 32668
rect 11472 32608 11536 32612
rect 14659 32668 14723 32672
rect 14659 32612 14663 32668
rect 14663 32612 14719 32668
rect 14719 32612 14723 32668
rect 14659 32608 14723 32612
rect 14739 32668 14803 32672
rect 14739 32612 14743 32668
rect 14743 32612 14799 32668
rect 14799 32612 14803 32668
rect 14739 32608 14803 32612
rect 14819 32668 14883 32672
rect 14819 32612 14823 32668
rect 14823 32612 14879 32668
rect 14879 32612 14883 32668
rect 14819 32608 14883 32612
rect 14899 32668 14963 32672
rect 14899 32612 14903 32668
rect 14903 32612 14959 32668
rect 14959 32612 14963 32668
rect 14899 32608 14963 32612
rect 2665 32124 2729 32128
rect 2665 32068 2669 32124
rect 2669 32068 2725 32124
rect 2725 32068 2729 32124
rect 2665 32064 2729 32068
rect 2745 32124 2809 32128
rect 2745 32068 2749 32124
rect 2749 32068 2805 32124
rect 2805 32068 2809 32124
rect 2745 32064 2809 32068
rect 2825 32124 2889 32128
rect 2825 32068 2829 32124
rect 2829 32068 2885 32124
rect 2885 32068 2889 32124
rect 2825 32064 2889 32068
rect 2905 32124 2969 32128
rect 2905 32068 2909 32124
rect 2909 32068 2965 32124
rect 2965 32068 2969 32124
rect 2905 32064 2969 32068
rect 6092 32124 6156 32128
rect 6092 32068 6096 32124
rect 6096 32068 6152 32124
rect 6152 32068 6156 32124
rect 6092 32064 6156 32068
rect 6172 32124 6236 32128
rect 6172 32068 6176 32124
rect 6176 32068 6232 32124
rect 6232 32068 6236 32124
rect 6172 32064 6236 32068
rect 6252 32124 6316 32128
rect 6252 32068 6256 32124
rect 6256 32068 6312 32124
rect 6312 32068 6316 32124
rect 6252 32064 6316 32068
rect 6332 32124 6396 32128
rect 6332 32068 6336 32124
rect 6336 32068 6392 32124
rect 6392 32068 6396 32124
rect 6332 32064 6396 32068
rect 9519 32124 9583 32128
rect 9519 32068 9523 32124
rect 9523 32068 9579 32124
rect 9579 32068 9583 32124
rect 9519 32064 9583 32068
rect 9599 32124 9663 32128
rect 9599 32068 9603 32124
rect 9603 32068 9659 32124
rect 9659 32068 9663 32124
rect 9599 32064 9663 32068
rect 9679 32124 9743 32128
rect 9679 32068 9683 32124
rect 9683 32068 9739 32124
rect 9739 32068 9743 32124
rect 9679 32064 9743 32068
rect 9759 32124 9823 32128
rect 9759 32068 9763 32124
rect 9763 32068 9819 32124
rect 9819 32068 9823 32124
rect 9759 32064 9823 32068
rect 12946 32124 13010 32128
rect 12946 32068 12950 32124
rect 12950 32068 13006 32124
rect 13006 32068 13010 32124
rect 12946 32064 13010 32068
rect 13026 32124 13090 32128
rect 13026 32068 13030 32124
rect 13030 32068 13086 32124
rect 13086 32068 13090 32124
rect 13026 32064 13090 32068
rect 13106 32124 13170 32128
rect 13106 32068 13110 32124
rect 13110 32068 13166 32124
rect 13166 32068 13170 32124
rect 13106 32064 13170 32068
rect 13186 32124 13250 32128
rect 13186 32068 13190 32124
rect 13190 32068 13246 32124
rect 13246 32068 13250 32124
rect 13186 32064 13250 32068
rect 4378 31580 4442 31584
rect 4378 31524 4382 31580
rect 4382 31524 4438 31580
rect 4438 31524 4442 31580
rect 4378 31520 4442 31524
rect 4458 31580 4522 31584
rect 4458 31524 4462 31580
rect 4462 31524 4518 31580
rect 4518 31524 4522 31580
rect 4458 31520 4522 31524
rect 4538 31580 4602 31584
rect 4538 31524 4542 31580
rect 4542 31524 4598 31580
rect 4598 31524 4602 31580
rect 4538 31520 4602 31524
rect 4618 31580 4682 31584
rect 4618 31524 4622 31580
rect 4622 31524 4678 31580
rect 4678 31524 4682 31580
rect 4618 31520 4682 31524
rect 7805 31580 7869 31584
rect 7805 31524 7809 31580
rect 7809 31524 7865 31580
rect 7865 31524 7869 31580
rect 7805 31520 7869 31524
rect 7885 31580 7949 31584
rect 7885 31524 7889 31580
rect 7889 31524 7945 31580
rect 7945 31524 7949 31580
rect 7885 31520 7949 31524
rect 7965 31580 8029 31584
rect 7965 31524 7969 31580
rect 7969 31524 8025 31580
rect 8025 31524 8029 31580
rect 7965 31520 8029 31524
rect 8045 31580 8109 31584
rect 8045 31524 8049 31580
rect 8049 31524 8105 31580
rect 8105 31524 8109 31580
rect 8045 31520 8109 31524
rect 11232 31580 11296 31584
rect 11232 31524 11236 31580
rect 11236 31524 11292 31580
rect 11292 31524 11296 31580
rect 11232 31520 11296 31524
rect 11312 31580 11376 31584
rect 11312 31524 11316 31580
rect 11316 31524 11372 31580
rect 11372 31524 11376 31580
rect 11312 31520 11376 31524
rect 11392 31580 11456 31584
rect 11392 31524 11396 31580
rect 11396 31524 11452 31580
rect 11452 31524 11456 31580
rect 11392 31520 11456 31524
rect 11472 31580 11536 31584
rect 11472 31524 11476 31580
rect 11476 31524 11532 31580
rect 11532 31524 11536 31580
rect 11472 31520 11536 31524
rect 14659 31580 14723 31584
rect 14659 31524 14663 31580
rect 14663 31524 14719 31580
rect 14719 31524 14723 31580
rect 14659 31520 14723 31524
rect 14739 31580 14803 31584
rect 14739 31524 14743 31580
rect 14743 31524 14799 31580
rect 14799 31524 14803 31580
rect 14739 31520 14803 31524
rect 14819 31580 14883 31584
rect 14819 31524 14823 31580
rect 14823 31524 14879 31580
rect 14879 31524 14883 31580
rect 14819 31520 14883 31524
rect 14899 31580 14963 31584
rect 14899 31524 14903 31580
rect 14903 31524 14959 31580
rect 14959 31524 14963 31580
rect 14899 31520 14963 31524
rect 2665 31036 2729 31040
rect 2665 30980 2669 31036
rect 2669 30980 2725 31036
rect 2725 30980 2729 31036
rect 2665 30976 2729 30980
rect 2745 31036 2809 31040
rect 2745 30980 2749 31036
rect 2749 30980 2805 31036
rect 2805 30980 2809 31036
rect 2745 30976 2809 30980
rect 2825 31036 2889 31040
rect 2825 30980 2829 31036
rect 2829 30980 2885 31036
rect 2885 30980 2889 31036
rect 2825 30976 2889 30980
rect 2905 31036 2969 31040
rect 2905 30980 2909 31036
rect 2909 30980 2965 31036
rect 2965 30980 2969 31036
rect 2905 30976 2969 30980
rect 6092 31036 6156 31040
rect 6092 30980 6096 31036
rect 6096 30980 6152 31036
rect 6152 30980 6156 31036
rect 6092 30976 6156 30980
rect 6172 31036 6236 31040
rect 6172 30980 6176 31036
rect 6176 30980 6232 31036
rect 6232 30980 6236 31036
rect 6172 30976 6236 30980
rect 6252 31036 6316 31040
rect 6252 30980 6256 31036
rect 6256 30980 6312 31036
rect 6312 30980 6316 31036
rect 6252 30976 6316 30980
rect 6332 31036 6396 31040
rect 6332 30980 6336 31036
rect 6336 30980 6392 31036
rect 6392 30980 6396 31036
rect 6332 30976 6396 30980
rect 9519 31036 9583 31040
rect 9519 30980 9523 31036
rect 9523 30980 9579 31036
rect 9579 30980 9583 31036
rect 9519 30976 9583 30980
rect 9599 31036 9663 31040
rect 9599 30980 9603 31036
rect 9603 30980 9659 31036
rect 9659 30980 9663 31036
rect 9599 30976 9663 30980
rect 9679 31036 9743 31040
rect 9679 30980 9683 31036
rect 9683 30980 9739 31036
rect 9739 30980 9743 31036
rect 9679 30976 9743 30980
rect 9759 31036 9823 31040
rect 9759 30980 9763 31036
rect 9763 30980 9819 31036
rect 9819 30980 9823 31036
rect 9759 30976 9823 30980
rect 12946 31036 13010 31040
rect 12946 30980 12950 31036
rect 12950 30980 13006 31036
rect 13006 30980 13010 31036
rect 12946 30976 13010 30980
rect 13026 31036 13090 31040
rect 13026 30980 13030 31036
rect 13030 30980 13086 31036
rect 13086 30980 13090 31036
rect 13026 30976 13090 30980
rect 13106 31036 13170 31040
rect 13106 30980 13110 31036
rect 13110 30980 13166 31036
rect 13166 30980 13170 31036
rect 13106 30976 13170 30980
rect 13186 31036 13250 31040
rect 13186 30980 13190 31036
rect 13190 30980 13246 31036
rect 13246 30980 13250 31036
rect 13186 30976 13250 30980
rect 4378 30492 4442 30496
rect 4378 30436 4382 30492
rect 4382 30436 4438 30492
rect 4438 30436 4442 30492
rect 4378 30432 4442 30436
rect 4458 30492 4522 30496
rect 4458 30436 4462 30492
rect 4462 30436 4518 30492
rect 4518 30436 4522 30492
rect 4458 30432 4522 30436
rect 4538 30492 4602 30496
rect 4538 30436 4542 30492
rect 4542 30436 4598 30492
rect 4598 30436 4602 30492
rect 4538 30432 4602 30436
rect 4618 30492 4682 30496
rect 4618 30436 4622 30492
rect 4622 30436 4678 30492
rect 4678 30436 4682 30492
rect 4618 30432 4682 30436
rect 7805 30492 7869 30496
rect 7805 30436 7809 30492
rect 7809 30436 7865 30492
rect 7865 30436 7869 30492
rect 7805 30432 7869 30436
rect 7885 30492 7949 30496
rect 7885 30436 7889 30492
rect 7889 30436 7945 30492
rect 7945 30436 7949 30492
rect 7885 30432 7949 30436
rect 7965 30492 8029 30496
rect 7965 30436 7969 30492
rect 7969 30436 8025 30492
rect 8025 30436 8029 30492
rect 7965 30432 8029 30436
rect 8045 30492 8109 30496
rect 8045 30436 8049 30492
rect 8049 30436 8105 30492
rect 8105 30436 8109 30492
rect 8045 30432 8109 30436
rect 11232 30492 11296 30496
rect 11232 30436 11236 30492
rect 11236 30436 11292 30492
rect 11292 30436 11296 30492
rect 11232 30432 11296 30436
rect 11312 30492 11376 30496
rect 11312 30436 11316 30492
rect 11316 30436 11372 30492
rect 11372 30436 11376 30492
rect 11312 30432 11376 30436
rect 11392 30492 11456 30496
rect 11392 30436 11396 30492
rect 11396 30436 11452 30492
rect 11452 30436 11456 30492
rect 11392 30432 11456 30436
rect 11472 30492 11536 30496
rect 11472 30436 11476 30492
rect 11476 30436 11532 30492
rect 11532 30436 11536 30492
rect 11472 30432 11536 30436
rect 14659 30492 14723 30496
rect 14659 30436 14663 30492
rect 14663 30436 14719 30492
rect 14719 30436 14723 30492
rect 14659 30432 14723 30436
rect 14739 30492 14803 30496
rect 14739 30436 14743 30492
rect 14743 30436 14799 30492
rect 14799 30436 14803 30492
rect 14739 30432 14803 30436
rect 14819 30492 14883 30496
rect 14819 30436 14823 30492
rect 14823 30436 14879 30492
rect 14879 30436 14883 30492
rect 14819 30432 14883 30436
rect 14899 30492 14963 30496
rect 14899 30436 14903 30492
rect 14903 30436 14959 30492
rect 14959 30436 14963 30492
rect 14899 30432 14963 30436
rect 2665 29948 2729 29952
rect 2665 29892 2669 29948
rect 2669 29892 2725 29948
rect 2725 29892 2729 29948
rect 2665 29888 2729 29892
rect 2745 29948 2809 29952
rect 2745 29892 2749 29948
rect 2749 29892 2805 29948
rect 2805 29892 2809 29948
rect 2745 29888 2809 29892
rect 2825 29948 2889 29952
rect 2825 29892 2829 29948
rect 2829 29892 2885 29948
rect 2885 29892 2889 29948
rect 2825 29888 2889 29892
rect 2905 29948 2969 29952
rect 2905 29892 2909 29948
rect 2909 29892 2965 29948
rect 2965 29892 2969 29948
rect 2905 29888 2969 29892
rect 6092 29948 6156 29952
rect 6092 29892 6096 29948
rect 6096 29892 6152 29948
rect 6152 29892 6156 29948
rect 6092 29888 6156 29892
rect 6172 29948 6236 29952
rect 6172 29892 6176 29948
rect 6176 29892 6232 29948
rect 6232 29892 6236 29948
rect 6172 29888 6236 29892
rect 6252 29948 6316 29952
rect 6252 29892 6256 29948
rect 6256 29892 6312 29948
rect 6312 29892 6316 29948
rect 6252 29888 6316 29892
rect 6332 29948 6396 29952
rect 6332 29892 6336 29948
rect 6336 29892 6392 29948
rect 6392 29892 6396 29948
rect 6332 29888 6396 29892
rect 9519 29948 9583 29952
rect 9519 29892 9523 29948
rect 9523 29892 9579 29948
rect 9579 29892 9583 29948
rect 9519 29888 9583 29892
rect 9599 29948 9663 29952
rect 9599 29892 9603 29948
rect 9603 29892 9659 29948
rect 9659 29892 9663 29948
rect 9599 29888 9663 29892
rect 9679 29948 9743 29952
rect 9679 29892 9683 29948
rect 9683 29892 9739 29948
rect 9739 29892 9743 29948
rect 9679 29888 9743 29892
rect 9759 29948 9823 29952
rect 9759 29892 9763 29948
rect 9763 29892 9819 29948
rect 9819 29892 9823 29948
rect 9759 29888 9823 29892
rect 12946 29948 13010 29952
rect 12946 29892 12950 29948
rect 12950 29892 13006 29948
rect 13006 29892 13010 29948
rect 12946 29888 13010 29892
rect 13026 29948 13090 29952
rect 13026 29892 13030 29948
rect 13030 29892 13086 29948
rect 13086 29892 13090 29948
rect 13026 29888 13090 29892
rect 13106 29948 13170 29952
rect 13106 29892 13110 29948
rect 13110 29892 13166 29948
rect 13166 29892 13170 29948
rect 13106 29888 13170 29892
rect 13186 29948 13250 29952
rect 13186 29892 13190 29948
rect 13190 29892 13246 29948
rect 13246 29892 13250 29948
rect 13186 29888 13250 29892
rect 4378 29404 4442 29408
rect 4378 29348 4382 29404
rect 4382 29348 4438 29404
rect 4438 29348 4442 29404
rect 4378 29344 4442 29348
rect 4458 29404 4522 29408
rect 4458 29348 4462 29404
rect 4462 29348 4518 29404
rect 4518 29348 4522 29404
rect 4458 29344 4522 29348
rect 4538 29404 4602 29408
rect 4538 29348 4542 29404
rect 4542 29348 4598 29404
rect 4598 29348 4602 29404
rect 4538 29344 4602 29348
rect 4618 29404 4682 29408
rect 4618 29348 4622 29404
rect 4622 29348 4678 29404
rect 4678 29348 4682 29404
rect 4618 29344 4682 29348
rect 7805 29404 7869 29408
rect 7805 29348 7809 29404
rect 7809 29348 7865 29404
rect 7865 29348 7869 29404
rect 7805 29344 7869 29348
rect 7885 29404 7949 29408
rect 7885 29348 7889 29404
rect 7889 29348 7945 29404
rect 7945 29348 7949 29404
rect 7885 29344 7949 29348
rect 7965 29404 8029 29408
rect 7965 29348 7969 29404
rect 7969 29348 8025 29404
rect 8025 29348 8029 29404
rect 7965 29344 8029 29348
rect 8045 29404 8109 29408
rect 8045 29348 8049 29404
rect 8049 29348 8105 29404
rect 8105 29348 8109 29404
rect 8045 29344 8109 29348
rect 11232 29404 11296 29408
rect 11232 29348 11236 29404
rect 11236 29348 11292 29404
rect 11292 29348 11296 29404
rect 11232 29344 11296 29348
rect 11312 29404 11376 29408
rect 11312 29348 11316 29404
rect 11316 29348 11372 29404
rect 11372 29348 11376 29404
rect 11312 29344 11376 29348
rect 11392 29404 11456 29408
rect 11392 29348 11396 29404
rect 11396 29348 11452 29404
rect 11452 29348 11456 29404
rect 11392 29344 11456 29348
rect 11472 29404 11536 29408
rect 11472 29348 11476 29404
rect 11476 29348 11532 29404
rect 11532 29348 11536 29404
rect 11472 29344 11536 29348
rect 14659 29404 14723 29408
rect 14659 29348 14663 29404
rect 14663 29348 14719 29404
rect 14719 29348 14723 29404
rect 14659 29344 14723 29348
rect 14739 29404 14803 29408
rect 14739 29348 14743 29404
rect 14743 29348 14799 29404
rect 14799 29348 14803 29404
rect 14739 29344 14803 29348
rect 14819 29404 14883 29408
rect 14819 29348 14823 29404
rect 14823 29348 14879 29404
rect 14879 29348 14883 29404
rect 14819 29344 14883 29348
rect 14899 29404 14963 29408
rect 14899 29348 14903 29404
rect 14903 29348 14959 29404
rect 14959 29348 14963 29404
rect 14899 29344 14963 29348
rect 2665 28860 2729 28864
rect 2665 28804 2669 28860
rect 2669 28804 2725 28860
rect 2725 28804 2729 28860
rect 2665 28800 2729 28804
rect 2745 28860 2809 28864
rect 2745 28804 2749 28860
rect 2749 28804 2805 28860
rect 2805 28804 2809 28860
rect 2745 28800 2809 28804
rect 2825 28860 2889 28864
rect 2825 28804 2829 28860
rect 2829 28804 2885 28860
rect 2885 28804 2889 28860
rect 2825 28800 2889 28804
rect 2905 28860 2969 28864
rect 2905 28804 2909 28860
rect 2909 28804 2965 28860
rect 2965 28804 2969 28860
rect 2905 28800 2969 28804
rect 6092 28860 6156 28864
rect 6092 28804 6096 28860
rect 6096 28804 6152 28860
rect 6152 28804 6156 28860
rect 6092 28800 6156 28804
rect 6172 28860 6236 28864
rect 6172 28804 6176 28860
rect 6176 28804 6232 28860
rect 6232 28804 6236 28860
rect 6172 28800 6236 28804
rect 6252 28860 6316 28864
rect 6252 28804 6256 28860
rect 6256 28804 6312 28860
rect 6312 28804 6316 28860
rect 6252 28800 6316 28804
rect 6332 28860 6396 28864
rect 6332 28804 6336 28860
rect 6336 28804 6392 28860
rect 6392 28804 6396 28860
rect 6332 28800 6396 28804
rect 9519 28860 9583 28864
rect 9519 28804 9523 28860
rect 9523 28804 9579 28860
rect 9579 28804 9583 28860
rect 9519 28800 9583 28804
rect 9599 28860 9663 28864
rect 9599 28804 9603 28860
rect 9603 28804 9659 28860
rect 9659 28804 9663 28860
rect 9599 28800 9663 28804
rect 9679 28860 9743 28864
rect 9679 28804 9683 28860
rect 9683 28804 9739 28860
rect 9739 28804 9743 28860
rect 9679 28800 9743 28804
rect 9759 28860 9823 28864
rect 9759 28804 9763 28860
rect 9763 28804 9819 28860
rect 9819 28804 9823 28860
rect 9759 28800 9823 28804
rect 12946 28860 13010 28864
rect 12946 28804 12950 28860
rect 12950 28804 13006 28860
rect 13006 28804 13010 28860
rect 12946 28800 13010 28804
rect 13026 28860 13090 28864
rect 13026 28804 13030 28860
rect 13030 28804 13086 28860
rect 13086 28804 13090 28860
rect 13026 28800 13090 28804
rect 13106 28860 13170 28864
rect 13106 28804 13110 28860
rect 13110 28804 13166 28860
rect 13166 28804 13170 28860
rect 13106 28800 13170 28804
rect 13186 28860 13250 28864
rect 13186 28804 13190 28860
rect 13190 28804 13246 28860
rect 13246 28804 13250 28860
rect 13186 28800 13250 28804
rect 4378 28316 4442 28320
rect 4378 28260 4382 28316
rect 4382 28260 4438 28316
rect 4438 28260 4442 28316
rect 4378 28256 4442 28260
rect 4458 28316 4522 28320
rect 4458 28260 4462 28316
rect 4462 28260 4518 28316
rect 4518 28260 4522 28316
rect 4458 28256 4522 28260
rect 4538 28316 4602 28320
rect 4538 28260 4542 28316
rect 4542 28260 4598 28316
rect 4598 28260 4602 28316
rect 4538 28256 4602 28260
rect 4618 28316 4682 28320
rect 4618 28260 4622 28316
rect 4622 28260 4678 28316
rect 4678 28260 4682 28316
rect 4618 28256 4682 28260
rect 7805 28316 7869 28320
rect 7805 28260 7809 28316
rect 7809 28260 7865 28316
rect 7865 28260 7869 28316
rect 7805 28256 7869 28260
rect 7885 28316 7949 28320
rect 7885 28260 7889 28316
rect 7889 28260 7945 28316
rect 7945 28260 7949 28316
rect 7885 28256 7949 28260
rect 7965 28316 8029 28320
rect 7965 28260 7969 28316
rect 7969 28260 8025 28316
rect 8025 28260 8029 28316
rect 7965 28256 8029 28260
rect 8045 28316 8109 28320
rect 8045 28260 8049 28316
rect 8049 28260 8105 28316
rect 8105 28260 8109 28316
rect 8045 28256 8109 28260
rect 11232 28316 11296 28320
rect 11232 28260 11236 28316
rect 11236 28260 11292 28316
rect 11292 28260 11296 28316
rect 11232 28256 11296 28260
rect 11312 28316 11376 28320
rect 11312 28260 11316 28316
rect 11316 28260 11372 28316
rect 11372 28260 11376 28316
rect 11312 28256 11376 28260
rect 11392 28316 11456 28320
rect 11392 28260 11396 28316
rect 11396 28260 11452 28316
rect 11452 28260 11456 28316
rect 11392 28256 11456 28260
rect 11472 28316 11536 28320
rect 11472 28260 11476 28316
rect 11476 28260 11532 28316
rect 11532 28260 11536 28316
rect 11472 28256 11536 28260
rect 14659 28316 14723 28320
rect 14659 28260 14663 28316
rect 14663 28260 14719 28316
rect 14719 28260 14723 28316
rect 14659 28256 14723 28260
rect 14739 28316 14803 28320
rect 14739 28260 14743 28316
rect 14743 28260 14799 28316
rect 14799 28260 14803 28316
rect 14739 28256 14803 28260
rect 14819 28316 14883 28320
rect 14819 28260 14823 28316
rect 14823 28260 14879 28316
rect 14879 28260 14883 28316
rect 14819 28256 14883 28260
rect 14899 28316 14963 28320
rect 14899 28260 14903 28316
rect 14903 28260 14959 28316
rect 14959 28260 14963 28316
rect 14899 28256 14963 28260
rect 2665 27772 2729 27776
rect 2665 27716 2669 27772
rect 2669 27716 2725 27772
rect 2725 27716 2729 27772
rect 2665 27712 2729 27716
rect 2745 27772 2809 27776
rect 2745 27716 2749 27772
rect 2749 27716 2805 27772
rect 2805 27716 2809 27772
rect 2745 27712 2809 27716
rect 2825 27772 2889 27776
rect 2825 27716 2829 27772
rect 2829 27716 2885 27772
rect 2885 27716 2889 27772
rect 2825 27712 2889 27716
rect 2905 27772 2969 27776
rect 2905 27716 2909 27772
rect 2909 27716 2965 27772
rect 2965 27716 2969 27772
rect 2905 27712 2969 27716
rect 6092 27772 6156 27776
rect 6092 27716 6096 27772
rect 6096 27716 6152 27772
rect 6152 27716 6156 27772
rect 6092 27712 6156 27716
rect 6172 27772 6236 27776
rect 6172 27716 6176 27772
rect 6176 27716 6232 27772
rect 6232 27716 6236 27772
rect 6172 27712 6236 27716
rect 6252 27772 6316 27776
rect 6252 27716 6256 27772
rect 6256 27716 6312 27772
rect 6312 27716 6316 27772
rect 6252 27712 6316 27716
rect 6332 27772 6396 27776
rect 6332 27716 6336 27772
rect 6336 27716 6392 27772
rect 6392 27716 6396 27772
rect 6332 27712 6396 27716
rect 9519 27772 9583 27776
rect 9519 27716 9523 27772
rect 9523 27716 9579 27772
rect 9579 27716 9583 27772
rect 9519 27712 9583 27716
rect 9599 27772 9663 27776
rect 9599 27716 9603 27772
rect 9603 27716 9659 27772
rect 9659 27716 9663 27772
rect 9599 27712 9663 27716
rect 9679 27772 9743 27776
rect 9679 27716 9683 27772
rect 9683 27716 9739 27772
rect 9739 27716 9743 27772
rect 9679 27712 9743 27716
rect 9759 27772 9823 27776
rect 9759 27716 9763 27772
rect 9763 27716 9819 27772
rect 9819 27716 9823 27772
rect 9759 27712 9823 27716
rect 12946 27772 13010 27776
rect 12946 27716 12950 27772
rect 12950 27716 13006 27772
rect 13006 27716 13010 27772
rect 12946 27712 13010 27716
rect 13026 27772 13090 27776
rect 13026 27716 13030 27772
rect 13030 27716 13086 27772
rect 13086 27716 13090 27772
rect 13026 27712 13090 27716
rect 13106 27772 13170 27776
rect 13106 27716 13110 27772
rect 13110 27716 13166 27772
rect 13166 27716 13170 27772
rect 13106 27712 13170 27716
rect 13186 27772 13250 27776
rect 13186 27716 13190 27772
rect 13190 27716 13246 27772
rect 13246 27716 13250 27772
rect 13186 27712 13250 27716
rect 4378 27228 4442 27232
rect 4378 27172 4382 27228
rect 4382 27172 4438 27228
rect 4438 27172 4442 27228
rect 4378 27168 4442 27172
rect 4458 27228 4522 27232
rect 4458 27172 4462 27228
rect 4462 27172 4518 27228
rect 4518 27172 4522 27228
rect 4458 27168 4522 27172
rect 4538 27228 4602 27232
rect 4538 27172 4542 27228
rect 4542 27172 4598 27228
rect 4598 27172 4602 27228
rect 4538 27168 4602 27172
rect 4618 27228 4682 27232
rect 4618 27172 4622 27228
rect 4622 27172 4678 27228
rect 4678 27172 4682 27228
rect 4618 27168 4682 27172
rect 7805 27228 7869 27232
rect 7805 27172 7809 27228
rect 7809 27172 7865 27228
rect 7865 27172 7869 27228
rect 7805 27168 7869 27172
rect 7885 27228 7949 27232
rect 7885 27172 7889 27228
rect 7889 27172 7945 27228
rect 7945 27172 7949 27228
rect 7885 27168 7949 27172
rect 7965 27228 8029 27232
rect 7965 27172 7969 27228
rect 7969 27172 8025 27228
rect 8025 27172 8029 27228
rect 7965 27168 8029 27172
rect 8045 27228 8109 27232
rect 8045 27172 8049 27228
rect 8049 27172 8105 27228
rect 8105 27172 8109 27228
rect 8045 27168 8109 27172
rect 11232 27228 11296 27232
rect 11232 27172 11236 27228
rect 11236 27172 11292 27228
rect 11292 27172 11296 27228
rect 11232 27168 11296 27172
rect 11312 27228 11376 27232
rect 11312 27172 11316 27228
rect 11316 27172 11372 27228
rect 11372 27172 11376 27228
rect 11312 27168 11376 27172
rect 11392 27228 11456 27232
rect 11392 27172 11396 27228
rect 11396 27172 11452 27228
rect 11452 27172 11456 27228
rect 11392 27168 11456 27172
rect 11472 27228 11536 27232
rect 11472 27172 11476 27228
rect 11476 27172 11532 27228
rect 11532 27172 11536 27228
rect 11472 27168 11536 27172
rect 14659 27228 14723 27232
rect 14659 27172 14663 27228
rect 14663 27172 14719 27228
rect 14719 27172 14723 27228
rect 14659 27168 14723 27172
rect 14739 27228 14803 27232
rect 14739 27172 14743 27228
rect 14743 27172 14799 27228
rect 14799 27172 14803 27228
rect 14739 27168 14803 27172
rect 14819 27228 14883 27232
rect 14819 27172 14823 27228
rect 14823 27172 14879 27228
rect 14879 27172 14883 27228
rect 14819 27168 14883 27172
rect 14899 27228 14963 27232
rect 14899 27172 14903 27228
rect 14903 27172 14959 27228
rect 14959 27172 14963 27228
rect 14899 27168 14963 27172
rect 2665 26684 2729 26688
rect 2665 26628 2669 26684
rect 2669 26628 2725 26684
rect 2725 26628 2729 26684
rect 2665 26624 2729 26628
rect 2745 26684 2809 26688
rect 2745 26628 2749 26684
rect 2749 26628 2805 26684
rect 2805 26628 2809 26684
rect 2745 26624 2809 26628
rect 2825 26684 2889 26688
rect 2825 26628 2829 26684
rect 2829 26628 2885 26684
rect 2885 26628 2889 26684
rect 2825 26624 2889 26628
rect 2905 26684 2969 26688
rect 2905 26628 2909 26684
rect 2909 26628 2965 26684
rect 2965 26628 2969 26684
rect 2905 26624 2969 26628
rect 6092 26684 6156 26688
rect 6092 26628 6096 26684
rect 6096 26628 6152 26684
rect 6152 26628 6156 26684
rect 6092 26624 6156 26628
rect 6172 26684 6236 26688
rect 6172 26628 6176 26684
rect 6176 26628 6232 26684
rect 6232 26628 6236 26684
rect 6172 26624 6236 26628
rect 6252 26684 6316 26688
rect 6252 26628 6256 26684
rect 6256 26628 6312 26684
rect 6312 26628 6316 26684
rect 6252 26624 6316 26628
rect 6332 26684 6396 26688
rect 6332 26628 6336 26684
rect 6336 26628 6392 26684
rect 6392 26628 6396 26684
rect 6332 26624 6396 26628
rect 9519 26684 9583 26688
rect 9519 26628 9523 26684
rect 9523 26628 9579 26684
rect 9579 26628 9583 26684
rect 9519 26624 9583 26628
rect 9599 26684 9663 26688
rect 9599 26628 9603 26684
rect 9603 26628 9659 26684
rect 9659 26628 9663 26684
rect 9599 26624 9663 26628
rect 9679 26684 9743 26688
rect 9679 26628 9683 26684
rect 9683 26628 9739 26684
rect 9739 26628 9743 26684
rect 9679 26624 9743 26628
rect 9759 26684 9823 26688
rect 9759 26628 9763 26684
rect 9763 26628 9819 26684
rect 9819 26628 9823 26684
rect 9759 26624 9823 26628
rect 12946 26684 13010 26688
rect 12946 26628 12950 26684
rect 12950 26628 13006 26684
rect 13006 26628 13010 26684
rect 12946 26624 13010 26628
rect 13026 26684 13090 26688
rect 13026 26628 13030 26684
rect 13030 26628 13086 26684
rect 13086 26628 13090 26684
rect 13026 26624 13090 26628
rect 13106 26684 13170 26688
rect 13106 26628 13110 26684
rect 13110 26628 13166 26684
rect 13166 26628 13170 26684
rect 13106 26624 13170 26628
rect 13186 26684 13250 26688
rect 13186 26628 13190 26684
rect 13190 26628 13246 26684
rect 13246 26628 13250 26684
rect 13186 26624 13250 26628
rect 4378 26140 4442 26144
rect 4378 26084 4382 26140
rect 4382 26084 4438 26140
rect 4438 26084 4442 26140
rect 4378 26080 4442 26084
rect 4458 26140 4522 26144
rect 4458 26084 4462 26140
rect 4462 26084 4518 26140
rect 4518 26084 4522 26140
rect 4458 26080 4522 26084
rect 4538 26140 4602 26144
rect 4538 26084 4542 26140
rect 4542 26084 4598 26140
rect 4598 26084 4602 26140
rect 4538 26080 4602 26084
rect 4618 26140 4682 26144
rect 4618 26084 4622 26140
rect 4622 26084 4678 26140
rect 4678 26084 4682 26140
rect 4618 26080 4682 26084
rect 7805 26140 7869 26144
rect 7805 26084 7809 26140
rect 7809 26084 7865 26140
rect 7865 26084 7869 26140
rect 7805 26080 7869 26084
rect 7885 26140 7949 26144
rect 7885 26084 7889 26140
rect 7889 26084 7945 26140
rect 7945 26084 7949 26140
rect 7885 26080 7949 26084
rect 7965 26140 8029 26144
rect 7965 26084 7969 26140
rect 7969 26084 8025 26140
rect 8025 26084 8029 26140
rect 7965 26080 8029 26084
rect 8045 26140 8109 26144
rect 8045 26084 8049 26140
rect 8049 26084 8105 26140
rect 8105 26084 8109 26140
rect 8045 26080 8109 26084
rect 11232 26140 11296 26144
rect 11232 26084 11236 26140
rect 11236 26084 11292 26140
rect 11292 26084 11296 26140
rect 11232 26080 11296 26084
rect 11312 26140 11376 26144
rect 11312 26084 11316 26140
rect 11316 26084 11372 26140
rect 11372 26084 11376 26140
rect 11312 26080 11376 26084
rect 11392 26140 11456 26144
rect 11392 26084 11396 26140
rect 11396 26084 11452 26140
rect 11452 26084 11456 26140
rect 11392 26080 11456 26084
rect 11472 26140 11536 26144
rect 11472 26084 11476 26140
rect 11476 26084 11532 26140
rect 11532 26084 11536 26140
rect 11472 26080 11536 26084
rect 14659 26140 14723 26144
rect 14659 26084 14663 26140
rect 14663 26084 14719 26140
rect 14719 26084 14723 26140
rect 14659 26080 14723 26084
rect 14739 26140 14803 26144
rect 14739 26084 14743 26140
rect 14743 26084 14799 26140
rect 14799 26084 14803 26140
rect 14739 26080 14803 26084
rect 14819 26140 14883 26144
rect 14819 26084 14823 26140
rect 14823 26084 14879 26140
rect 14879 26084 14883 26140
rect 14819 26080 14883 26084
rect 14899 26140 14963 26144
rect 14899 26084 14903 26140
rect 14903 26084 14959 26140
rect 14959 26084 14963 26140
rect 14899 26080 14963 26084
rect 2665 25596 2729 25600
rect 2665 25540 2669 25596
rect 2669 25540 2725 25596
rect 2725 25540 2729 25596
rect 2665 25536 2729 25540
rect 2745 25596 2809 25600
rect 2745 25540 2749 25596
rect 2749 25540 2805 25596
rect 2805 25540 2809 25596
rect 2745 25536 2809 25540
rect 2825 25596 2889 25600
rect 2825 25540 2829 25596
rect 2829 25540 2885 25596
rect 2885 25540 2889 25596
rect 2825 25536 2889 25540
rect 2905 25596 2969 25600
rect 2905 25540 2909 25596
rect 2909 25540 2965 25596
rect 2965 25540 2969 25596
rect 2905 25536 2969 25540
rect 6092 25596 6156 25600
rect 6092 25540 6096 25596
rect 6096 25540 6152 25596
rect 6152 25540 6156 25596
rect 6092 25536 6156 25540
rect 6172 25596 6236 25600
rect 6172 25540 6176 25596
rect 6176 25540 6232 25596
rect 6232 25540 6236 25596
rect 6172 25536 6236 25540
rect 6252 25596 6316 25600
rect 6252 25540 6256 25596
rect 6256 25540 6312 25596
rect 6312 25540 6316 25596
rect 6252 25536 6316 25540
rect 6332 25596 6396 25600
rect 6332 25540 6336 25596
rect 6336 25540 6392 25596
rect 6392 25540 6396 25596
rect 6332 25536 6396 25540
rect 9519 25596 9583 25600
rect 9519 25540 9523 25596
rect 9523 25540 9579 25596
rect 9579 25540 9583 25596
rect 9519 25536 9583 25540
rect 9599 25596 9663 25600
rect 9599 25540 9603 25596
rect 9603 25540 9659 25596
rect 9659 25540 9663 25596
rect 9599 25536 9663 25540
rect 9679 25596 9743 25600
rect 9679 25540 9683 25596
rect 9683 25540 9739 25596
rect 9739 25540 9743 25596
rect 9679 25536 9743 25540
rect 9759 25596 9823 25600
rect 9759 25540 9763 25596
rect 9763 25540 9819 25596
rect 9819 25540 9823 25596
rect 9759 25536 9823 25540
rect 12946 25596 13010 25600
rect 12946 25540 12950 25596
rect 12950 25540 13006 25596
rect 13006 25540 13010 25596
rect 12946 25536 13010 25540
rect 13026 25596 13090 25600
rect 13026 25540 13030 25596
rect 13030 25540 13086 25596
rect 13086 25540 13090 25596
rect 13026 25536 13090 25540
rect 13106 25596 13170 25600
rect 13106 25540 13110 25596
rect 13110 25540 13166 25596
rect 13166 25540 13170 25596
rect 13106 25536 13170 25540
rect 13186 25596 13250 25600
rect 13186 25540 13190 25596
rect 13190 25540 13246 25596
rect 13246 25540 13250 25596
rect 13186 25536 13250 25540
rect 4378 25052 4442 25056
rect 4378 24996 4382 25052
rect 4382 24996 4438 25052
rect 4438 24996 4442 25052
rect 4378 24992 4442 24996
rect 4458 25052 4522 25056
rect 4458 24996 4462 25052
rect 4462 24996 4518 25052
rect 4518 24996 4522 25052
rect 4458 24992 4522 24996
rect 4538 25052 4602 25056
rect 4538 24996 4542 25052
rect 4542 24996 4598 25052
rect 4598 24996 4602 25052
rect 4538 24992 4602 24996
rect 4618 25052 4682 25056
rect 4618 24996 4622 25052
rect 4622 24996 4678 25052
rect 4678 24996 4682 25052
rect 4618 24992 4682 24996
rect 7805 25052 7869 25056
rect 7805 24996 7809 25052
rect 7809 24996 7865 25052
rect 7865 24996 7869 25052
rect 7805 24992 7869 24996
rect 7885 25052 7949 25056
rect 7885 24996 7889 25052
rect 7889 24996 7945 25052
rect 7945 24996 7949 25052
rect 7885 24992 7949 24996
rect 7965 25052 8029 25056
rect 7965 24996 7969 25052
rect 7969 24996 8025 25052
rect 8025 24996 8029 25052
rect 7965 24992 8029 24996
rect 8045 25052 8109 25056
rect 8045 24996 8049 25052
rect 8049 24996 8105 25052
rect 8105 24996 8109 25052
rect 8045 24992 8109 24996
rect 11232 25052 11296 25056
rect 11232 24996 11236 25052
rect 11236 24996 11292 25052
rect 11292 24996 11296 25052
rect 11232 24992 11296 24996
rect 11312 25052 11376 25056
rect 11312 24996 11316 25052
rect 11316 24996 11372 25052
rect 11372 24996 11376 25052
rect 11312 24992 11376 24996
rect 11392 25052 11456 25056
rect 11392 24996 11396 25052
rect 11396 24996 11452 25052
rect 11452 24996 11456 25052
rect 11392 24992 11456 24996
rect 11472 25052 11536 25056
rect 11472 24996 11476 25052
rect 11476 24996 11532 25052
rect 11532 24996 11536 25052
rect 11472 24992 11536 24996
rect 14659 25052 14723 25056
rect 14659 24996 14663 25052
rect 14663 24996 14719 25052
rect 14719 24996 14723 25052
rect 14659 24992 14723 24996
rect 14739 25052 14803 25056
rect 14739 24996 14743 25052
rect 14743 24996 14799 25052
rect 14799 24996 14803 25052
rect 14739 24992 14803 24996
rect 14819 25052 14883 25056
rect 14819 24996 14823 25052
rect 14823 24996 14879 25052
rect 14879 24996 14883 25052
rect 14819 24992 14883 24996
rect 14899 25052 14963 25056
rect 14899 24996 14903 25052
rect 14903 24996 14959 25052
rect 14959 24996 14963 25052
rect 14899 24992 14963 24996
rect 2665 24508 2729 24512
rect 2665 24452 2669 24508
rect 2669 24452 2725 24508
rect 2725 24452 2729 24508
rect 2665 24448 2729 24452
rect 2745 24508 2809 24512
rect 2745 24452 2749 24508
rect 2749 24452 2805 24508
rect 2805 24452 2809 24508
rect 2745 24448 2809 24452
rect 2825 24508 2889 24512
rect 2825 24452 2829 24508
rect 2829 24452 2885 24508
rect 2885 24452 2889 24508
rect 2825 24448 2889 24452
rect 2905 24508 2969 24512
rect 2905 24452 2909 24508
rect 2909 24452 2965 24508
rect 2965 24452 2969 24508
rect 2905 24448 2969 24452
rect 6092 24508 6156 24512
rect 6092 24452 6096 24508
rect 6096 24452 6152 24508
rect 6152 24452 6156 24508
rect 6092 24448 6156 24452
rect 6172 24508 6236 24512
rect 6172 24452 6176 24508
rect 6176 24452 6232 24508
rect 6232 24452 6236 24508
rect 6172 24448 6236 24452
rect 6252 24508 6316 24512
rect 6252 24452 6256 24508
rect 6256 24452 6312 24508
rect 6312 24452 6316 24508
rect 6252 24448 6316 24452
rect 6332 24508 6396 24512
rect 6332 24452 6336 24508
rect 6336 24452 6392 24508
rect 6392 24452 6396 24508
rect 6332 24448 6396 24452
rect 9519 24508 9583 24512
rect 9519 24452 9523 24508
rect 9523 24452 9579 24508
rect 9579 24452 9583 24508
rect 9519 24448 9583 24452
rect 9599 24508 9663 24512
rect 9599 24452 9603 24508
rect 9603 24452 9659 24508
rect 9659 24452 9663 24508
rect 9599 24448 9663 24452
rect 9679 24508 9743 24512
rect 9679 24452 9683 24508
rect 9683 24452 9739 24508
rect 9739 24452 9743 24508
rect 9679 24448 9743 24452
rect 9759 24508 9823 24512
rect 9759 24452 9763 24508
rect 9763 24452 9819 24508
rect 9819 24452 9823 24508
rect 9759 24448 9823 24452
rect 12946 24508 13010 24512
rect 12946 24452 12950 24508
rect 12950 24452 13006 24508
rect 13006 24452 13010 24508
rect 12946 24448 13010 24452
rect 13026 24508 13090 24512
rect 13026 24452 13030 24508
rect 13030 24452 13086 24508
rect 13086 24452 13090 24508
rect 13026 24448 13090 24452
rect 13106 24508 13170 24512
rect 13106 24452 13110 24508
rect 13110 24452 13166 24508
rect 13166 24452 13170 24508
rect 13106 24448 13170 24452
rect 13186 24508 13250 24512
rect 13186 24452 13190 24508
rect 13190 24452 13246 24508
rect 13246 24452 13250 24508
rect 13186 24448 13250 24452
rect 4378 23964 4442 23968
rect 4378 23908 4382 23964
rect 4382 23908 4438 23964
rect 4438 23908 4442 23964
rect 4378 23904 4442 23908
rect 4458 23964 4522 23968
rect 4458 23908 4462 23964
rect 4462 23908 4518 23964
rect 4518 23908 4522 23964
rect 4458 23904 4522 23908
rect 4538 23964 4602 23968
rect 4538 23908 4542 23964
rect 4542 23908 4598 23964
rect 4598 23908 4602 23964
rect 4538 23904 4602 23908
rect 4618 23964 4682 23968
rect 4618 23908 4622 23964
rect 4622 23908 4678 23964
rect 4678 23908 4682 23964
rect 4618 23904 4682 23908
rect 7805 23964 7869 23968
rect 7805 23908 7809 23964
rect 7809 23908 7865 23964
rect 7865 23908 7869 23964
rect 7805 23904 7869 23908
rect 7885 23964 7949 23968
rect 7885 23908 7889 23964
rect 7889 23908 7945 23964
rect 7945 23908 7949 23964
rect 7885 23904 7949 23908
rect 7965 23964 8029 23968
rect 7965 23908 7969 23964
rect 7969 23908 8025 23964
rect 8025 23908 8029 23964
rect 7965 23904 8029 23908
rect 8045 23964 8109 23968
rect 8045 23908 8049 23964
rect 8049 23908 8105 23964
rect 8105 23908 8109 23964
rect 8045 23904 8109 23908
rect 11232 23964 11296 23968
rect 11232 23908 11236 23964
rect 11236 23908 11292 23964
rect 11292 23908 11296 23964
rect 11232 23904 11296 23908
rect 11312 23964 11376 23968
rect 11312 23908 11316 23964
rect 11316 23908 11372 23964
rect 11372 23908 11376 23964
rect 11312 23904 11376 23908
rect 11392 23964 11456 23968
rect 11392 23908 11396 23964
rect 11396 23908 11452 23964
rect 11452 23908 11456 23964
rect 11392 23904 11456 23908
rect 11472 23964 11536 23968
rect 11472 23908 11476 23964
rect 11476 23908 11532 23964
rect 11532 23908 11536 23964
rect 11472 23904 11536 23908
rect 14659 23964 14723 23968
rect 14659 23908 14663 23964
rect 14663 23908 14719 23964
rect 14719 23908 14723 23964
rect 14659 23904 14723 23908
rect 14739 23964 14803 23968
rect 14739 23908 14743 23964
rect 14743 23908 14799 23964
rect 14799 23908 14803 23964
rect 14739 23904 14803 23908
rect 14819 23964 14883 23968
rect 14819 23908 14823 23964
rect 14823 23908 14879 23964
rect 14879 23908 14883 23964
rect 14819 23904 14883 23908
rect 14899 23964 14963 23968
rect 14899 23908 14903 23964
rect 14903 23908 14959 23964
rect 14959 23908 14963 23964
rect 14899 23904 14963 23908
rect 2665 23420 2729 23424
rect 2665 23364 2669 23420
rect 2669 23364 2725 23420
rect 2725 23364 2729 23420
rect 2665 23360 2729 23364
rect 2745 23420 2809 23424
rect 2745 23364 2749 23420
rect 2749 23364 2805 23420
rect 2805 23364 2809 23420
rect 2745 23360 2809 23364
rect 2825 23420 2889 23424
rect 2825 23364 2829 23420
rect 2829 23364 2885 23420
rect 2885 23364 2889 23420
rect 2825 23360 2889 23364
rect 2905 23420 2969 23424
rect 2905 23364 2909 23420
rect 2909 23364 2965 23420
rect 2965 23364 2969 23420
rect 2905 23360 2969 23364
rect 6092 23420 6156 23424
rect 6092 23364 6096 23420
rect 6096 23364 6152 23420
rect 6152 23364 6156 23420
rect 6092 23360 6156 23364
rect 6172 23420 6236 23424
rect 6172 23364 6176 23420
rect 6176 23364 6232 23420
rect 6232 23364 6236 23420
rect 6172 23360 6236 23364
rect 6252 23420 6316 23424
rect 6252 23364 6256 23420
rect 6256 23364 6312 23420
rect 6312 23364 6316 23420
rect 6252 23360 6316 23364
rect 6332 23420 6396 23424
rect 6332 23364 6336 23420
rect 6336 23364 6392 23420
rect 6392 23364 6396 23420
rect 6332 23360 6396 23364
rect 9519 23420 9583 23424
rect 9519 23364 9523 23420
rect 9523 23364 9579 23420
rect 9579 23364 9583 23420
rect 9519 23360 9583 23364
rect 9599 23420 9663 23424
rect 9599 23364 9603 23420
rect 9603 23364 9659 23420
rect 9659 23364 9663 23420
rect 9599 23360 9663 23364
rect 9679 23420 9743 23424
rect 9679 23364 9683 23420
rect 9683 23364 9739 23420
rect 9739 23364 9743 23420
rect 9679 23360 9743 23364
rect 9759 23420 9823 23424
rect 9759 23364 9763 23420
rect 9763 23364 9819 23420
rect 9819 23364 9823 23420
rect 9759 23360 9823 23364
rect 12946 23420 13010 23424
rect 12946 23364 12950 23420
rect 12950 23364 13006 23420
rect 13006 23364 13010 23420
rect 12946 23360 13010 23364
rect 13026 23420 13090 23424
rect 13026 23364 13030 23420
rect 13030 23364 13086 23420
rect 13086 23364 13090 23420
rect 13026 23360 13090 23364
rect 13106 23420 13170 23424
rect 13106 23364 13110 23420
rect 13110 23364 13166 23420
rect 13166 23364 13170 23420
rect 13106 23360 13170 23364
rect 13186 23420 13250 23424
rect 13186 23364 13190 23420
rect 13190 23364 13246 23420
rect 13246 23364 13250 23420
rect 13186 23360 13250 23364
rect 4378 22876 4442 22880
rect 4378 22820 4382 22876
rect 4382 22820 4438 22876
rect 4438 22820 4442 22876
rect 4378 22816 4442 22820
rect 4458 22876 4522 22880
rect 4458 22820 4462 22876
rect 4462 22820 4518 22876
rect 4518 22820 4522 22876
rect 4458 22816 4522 22820
rect 4538 22876 4602 22880
rect 4538 22820 4542 22876
rect 4542 22820 4598 22876
rect 4598 22820 4602 22876
rect 4538 22816 4602 22820
rect 4618 22876 4682 22880
rect 4618 22820 4622 22876
rect 4622 22820 4678 22876
rect 4678 22820 4682 22876
rect 4618 22816 4682 22820
rect 7805 22876 7869 22880
rect 7805 22820 7809 22876
rect 7809 22820 7865 22876
rect 7865 22820 7869 22876
rect 7805 22816 7869 22820
rect 7885 22876 7949 22880
rect 7885 22820 7889 22876
rect 7889 22820 7945 22876
rect 7945 22820 7949 22876
rect 7885 22816 7949 22820
rect 7965 22876 8029 22880
rect 7965 22820 7969 22876
rect 7969 22820 8025 22876
rect 8025 22820 8029 22876
rect 7965 22816 8029 22820
rect 8045 22876 8109 22880
rect 8045 22820 8049 22876
rect 8049 22820 8105 22876
rect 8105 22820 8109 22876
rect 8045 22816 8109 22820
rect 11232 22876 11296 22880
rect 11232 22820 11236 22876
rect 11236 22820 11292 22876
rect 11292 22820 11296 22876
rect 11232 22816 11296 22820
rect 11312 22876 11376 22880
rect 11312 22820 11316 22876
rect 11316 22820 11372 22876
rect 11372 22820 11376 22876
rect 11312 22816 11376 22820
rect 11392 22876 11456 22880
rect 11392 22820 11396 22876
rect 11396 22820 11452 22876
rect 11452 22820 11456 22876
rect 11392 22816 11456 22820
rect 11472 22876 11536 22880
rect 11472 22820 11476 22876
rect 11476 22820 11532 22876
rect 11532 22820 11536 22876
rect 11472 22816 11536 22820
rect 14659 22876 14723 22880
rect 14659 22820 14663 22876
rect 14663 22820 14719 22876
rect 14719 22820 14723 22876
rect 14659 22816 14723 22820
rect 14739 22876 14803 22880
rect 14739 22820 14743 22876
rect 14743 22820 14799 22876
rect 14799 22820 14803 22876
rect 14739 22816 14803 22820
rect 14819 22876 14883 22880
rect 14819 22820 14823 22876
rect 14823 22820 14879 22876
rect 14879 22820 14883 22876
rect 14819 22816 14883 22820
rect 14899 22876 14963 22880
rect 14899 22820 14903 22876
rect 14903 22820 14959 22876
rect 14959 22820 14963 22876
rect 14899 22816 14963 22820
rect 2665 22332 2729 22336
rect 2665 22276 2669 22332
rect 2669 22276 2725 22332
rect 2725 22276 2729 22332
rect 2665 22272 2729 22276
rect 2745 22332 2809 22336
rect 2745 22276 2749 22332
rect 2749 22276 2805 22332
rect 2805 22276 2809 22332
rect 2745 22272 2809 22276
rect 2825 22332 2889 22336
rect 2825 22276 2829 22332
rect 2829 22276 2885 22332
rect 2885 22276 2889 22332
rect 2825 22272 2889 22276
rect 2905 22332 2969 22336
rect 2905 22276 2909 22332
rect 2909 22276 2965 22332
rect 2965 22276 2969 22332
rect 2905 22272 2969 22276
rect 6092 22332 6156 22336
rect 6092 22276 6096 22332
rect 6096 22276 6152 22332
rect 6152 22276 6156 22332
rect 6092 22272 6156 22276
rect 6172 22332 6236 22336
rect 6172 22276 6176 22332
rect 6176 22276 6232 22332
rect 6232 22276 6236 22332
rect 6172 22272 6236 22276
rect 6252 22332 6316 22336
rect 6252 22276 6256 22332
rect 6256 22276 6312 22332
rect 6312 22276 6316 22332
rect 6252 22272 6316 22276
rect 6332 22332 6396 22336
rect 6332 22276 6336 22332
rect 6336 22276 6392 22332
rect 6392 22276 6396 22332
rect 6332 22272 6396 22276
rect 9519 22332 9583 22336
rect 9519 22276 9523 22332
rect 9523 22276 9579 22332
rect 9579 22276 9583 22332
rect 9519 22272 9583 22276
rect 9599 22332 9663 22336
rect 9599 22276 9603 22332
rect 9603 22276 9659 22332
rect 9659 22276 9663 22332
rect 9599 22272 9663 22276
rect 9679 22332 9743 22336
rect 9679 22276 9683 22332
rect 9683 22276 9739 22332
rect 9739 22276 9743 22332
rect 9679 22272 9743 22276
rect 9759 22332 9823 22336
rect 9759 22276 9763 22332
rect 9763 22276 9819 22332
rect 9819 22276 9823 22332
rect 9759 22272 9823 22276
rect 12946 22332 13010 22336
rect 12946 22276 12950 22332
rect 12950 22276 13006 22332
rect 13006 22276 13010 22332
rect 12946 22272 13010 22276
rect 13026 22332 13090 22336
rect 13026 22276 13030 22332
rect 13030 22276 13086 22332
rect 13086 22276 13090 22332
rect 13026 22272 13090 22276
rect 13106 22332 13170 22336
rect 13106 22276 13110 22332
rect 13110 22276 13166 22332
rect 13166 22276 13170 22332
rect 13106 22272 13170 22276
rect 13186 22332 13250 22336
rect 13186 22276 13190 22332
rect 13190 22276 13246 22332
rect 13246 22276 13250 22332
rect 13186 22272 13250 22276
rect 4378 21788 4442 21792
rect 4378 21732 4382 21788
rect 4382 21732 4438 21788
rect 4438 21732 4442 21788
rect 4378 21728 4442 21732
rect 4458 21788 4522 21792
rect 4458 21732 4462 21788
rect 4462 21732 4518 21788
rect 4518 21732 4522 21788
rect 4458 21728 4522 21732
rect 4538 21788 4602 21792
rect 4538 21732 4542 21788
rect 4542 21732 4598 21788
rect 4598 21732 4602 21788
rect 4538 21728 4602 21732
rect 4618 21788 4682 21792
rect 4618 21732 4622 21788
rect 4622 21732 4678 21788
rect 4678 21732 4682 21788
rect 4618 21728 4682 21732
rect 7805 21788 7869 21792
rect 7805 21732 7809 21788
rect 7809 21732 7865 21788
rect 7865 21732 7869 21788
rect 7805 21728 7869 21732
rect 7885 21788 7949 21792
rect 7885 21732 7889 21788
rect 7889 21732 7945 21788
rect 7945 21732 7949 21788
rect 7885 21728 7949 21732
rect 7965 21788 8029 21792
rect 7965 21732 7969 21788
rect 7969 21732 8025 21788
rect 8025 21732 8029 21788
rect 7965 21728 8029 21732
rect 8045 21788 8109 21792
rect 8045 21732 8049 21788
rect 8049 21732 8105 21788
rect 8105 21732 8109 21788
rect 8045 21728 8109 21732
rect 11232 21788 11296 21792
rect 11232 21732 11236 21788
rect 11236 21732 11292 21788
rect 11292 21732 11296 21788
rect 11232 21728 11296 21732
rect 11312 21788 11376 21792
rect 11312 21732 11316 21788
rect 11316 21732 11372 21788
rect 11372 21732 11376 21788
rect 11312 21728 11376 21732
rect 11392 21788 11456 21792
rect 11392 21732 11396 21788
rect 11396 21732 11452 21788
rect 11452 21732 11456 21788
rect 11392 21728 11456 21732
rect 11472 21788 11536 21792
rect 11472 21732 11476 21788
rect 11476 21732 11532 21788
rect 11532 21732 11536 21788
rect 11472 21728 11536 21732
rect 14659 21788 14723 21792
rect 14659 21732 14663 21788
rect 14663 21732 14719 21788
rect 14719 21732 14723 21788
rect 14659 21728 14723 21732
rect 14739 21788 14803 21792
rect 14739 21732 14743 21788
rect 14743 21732 14799 21788
rect 14799 21732 14803 21788
rect 14739 21728 14803 21732
rect 14819 21788 14883 21792
rect 14819 21732 14823 21788
rect 14823 21732 14879 21788
rect 14879 21732 14883 21788
rect 14819 21728 14883 21732
rect 14899 21788 14963 21792
rect 14899 21732 14903 21788
rect 14903 21732 14959 21788
rect 14959 21732 14963 21788
rect 14899 21728 14963 21732
rect 2665 21244 2729 21248
rect 2665 21188 2669 21244
rect 2669 21188 2725 21244
rect 2725 21188 2729 21244
rect 2665 21184 2729 21188
rect 2745 21244 2809 21248
rect 2745 21188 2749 21244
rect 2749 21188 2805 21244
rect 2805 21188 2809 21244
rect 2745 21184 2809 21188
rect 2825 21244 2889 21248
rect 2825 21188 2829 21244
rect 2829 21188 2885 21244
rect 2885 21188 2889 21244
rect 2825 21184 2889 21188
rect 2905 21244 2969 21248
rect 2905 21188 2909 21244
rect 2909 21188 2965 21244
rect 2965 21188 2969 21244
rect 2905 21184 2969 21188
rect 6092 21244 6156 21248
rect 6092 21188 6096 21244
rect 6096 21188 6152 21244
rect 6152 21188 6156 21244
rect 6092 21184 6156 21188
rect 6172 21244 6236 21248
rect 6172 21188 6176 21244
rect 6176 21188 6232 21244
rect 6232 21188 6236 21244
rect 6172 21184 6236 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 9519 21244 9583 21248
rect 9519 21188 9523 21244
rect 9523 21188 9579 21244
rect 9579 21188 9583 21244
rect 9519 21184 9583 21188
rect 9599 21244 9663 21248
rect 9599 21188 9603 21244
rect 9603 21188 9659 21244
rect 9659 21188 9663 21244
rect 9599 21184 9663 21188
rect 9679 21244 9743 21248
rect 9679 21188 9683 21244
rect 9683 21188 9739 21244
rect 9739 21188 9743 21244
rect 9679 21184 9743 21188
rect 9759 21244 9823 21248
rect 9759 21188 9763 21244
rect 9763 21188 9819 21244
rect 9819 21188 9823 21244
rect 9759 21184 9823 21188
rect 12946 21244 13010 21248
rect 12946 21188 12950 21244
rect 12950 21188 13006 21244
rect 13006 21188 13010 21244
rect 12946 21184 13010 21188
rect 13026 21244 13090 21248
rect 13026 21188 13030 21244
rect 13030 21188 13086 21244
rect 13086 21188 13090 21244
rect 13026 21184 13090 21188
rect 13106 21244 13170 21248
rect 13106 21188 13110 21244
rect 13110 21188 13166 21244
rect 13166 21188 13170 21244
rect 13106 21184 13170 21188
rect 13186 21244 13250 21248
rect 13186 21188 13190 21244
rect 13190 21188 13246 21244
rect 13246 21188 13250 21244
rect 13186 21184 13250 21188
rect 4378 20700 4442 20704
rect 4378 20644 4382 20700
rect 4382 20644 4438 20700
rect 4438 20644 4442 20700
rect 4378 20640 4442 20644
rect 4458 20700 4522 20704
rect 4458 20644 4462 20700
rect 4462 20644 4518 20700
rect 4518 20644 4522 20700
rect 4458 20640 4522 20644
rect 4538 20700 4602 20704
rect 4538 20644 4542 20700
rect 4542 20644 4598 20700
rect 4598 20644 4602 20700
rect 4538 20640 4602 20644
rect 4618 20700 4682 20704
rect 4618 20644 4622 20700
rect 4622 20644 4678 20700
rect 4678 20644 4682 20700
rect 4618 20640 4682 20644
rect 7805 20700 7869 20704
rect 7805 20644 7809 20700
rect 7809 20644 7865 20700
rect 7865 20644 7869 20700
rect 7805 20640 7869 20644
rect 7885 20700 7949 20704
rect 7885 20644 7889 20700
rect 7889 20644 7945 20700
rect 7945 20644 7949 20700
rect 7885 20640 7949 20644
rect 7965 20700 8029 20704
rect 7965 20644 7969 20700
rect 7969 20644 8025 20700
rect 8025 20644 8029 20700
rect 7965 20640 8029 20644
rect 8045 20700 8109 20704
rect 8045 20644 8049 20700
rect 8049 20644 8105 20700
rect 8105 20644 8109 20700
rect 8045 20640 8109 20644
rect 11232 20700 11296 20704
rect 11232 20644 11236 20700
rect 11236 20644 11292 20700
rect 11292 20644 11296 20700
rect 11232 20640 11296 20644
rect 11312 20700 11376 20704
rect 11312 20644 11316 20700
rect 11316 20644 11372 20700
rect 11372 20644 11376 20700
rect 11312 20640 11376 20644
rect 11392 20700 11456 20704
rect 11392 20644 11396 20700
rect 11396 20644 11452 20700
rect 11452 20644 11456 20700
rect 11392 20640 11456 20644
rect 11472 20700 11536 20704
rect 11472 20644 11476 20700
rect 11476 20644 11532 20700
rect 11532 20644 11536 20700
rect 11472 20640 11536 20644
rect 14659 20700 14723 20704
rect 14659 20644 14663 20700
rect 14663 20644 14719 20700
rect 14719 20644 14723 20700
rect 14659 20640 14723 20644
rect 14739 20700 14803 20704
rect 14739 20644 14743 20700
rect 14743 20644 14799 20700
rect 14799 20644 14803 20700
rect 14739 20640 14803 20644
rect 14819 20700 14883 20704
rect 14819 20644 14823 20700
rect 14823 20644 14879 20700
rect 14879 20644 14883 20700
rect 14819 20640 14883 20644
rect 14899 20700 14963 20704
rect 14899 20644 14903 20700
rect 14903 20644 14959 20700
rect 14959 20644 14963 20700
rect 14899 20640 14963 20644
rect 2665 20156 2729 20160
rect 2665 20100 2669 20156
rect 2669 20100 2725 20156
rect 2725 20100 2729 20156
rect 2665 20096 2729 20100
rect 2745 20156 2809 20160
rect 2745 20100 2749 20156
rect 2749 20100 2805 20156
rect 2805 20100 2809 20156
rect 2745 20096 2809 20100
rect 2825 20156 2889 20160
rect 2825 20100 2829 20156
rect 2829 20100 2885 20156
rect 2885 20100 2889 20156
rect 2825 20096 2889 20100
rect 2905 20156 2969 20160
rect 2905 20100 2909 20156
rect 2909 20100 2965 20156
rect 2965 20100 2969 20156
rect 2905 20096 2969 20100
rect 6092 20156 6156 20160
rect 6092 20100 6096 20156
rect 6096 20100 6152 20156
rect 6152 20100 6156 20156
rect 6092 20096 6156 20100
rect 6172 20156 6236 20160
rect 6172 20100 6176 20156
rect 6176 20100 6232 20156
rect 6232 20100 6236 20156
rect 6172 20096 6236 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 9519 20156 9583 20160
rect 9519 20100 9523 20156
rect 9523 20100 9579 20156
rect 9579 20100 9583 20156
rect 9519 20096 9583 20100
rect 9599 20156 9663 20160
rect 9599 20100 9603 20156
rect 9603 20100 9659 20156
rect 9659 20100 9663 20156
rect 9599 20096 9663 20100
rect 9679 20156 9743 20160
rect 9679 20100 9683 20156
rect 9683 20100 9739 20156
rect 9739 20100 9743 20156
rect 9679 20096 9743 20100
rect 9759 20156 9823 20160
rect 9759 20100 9763 20156
rect 9763 20100 9819 20156
rect 9819 20100 9823 20156
rect 9759 20096 9823 20100
rect 12946 20156 13010 20160
rect 12946 20100 12950 20156
rect 12950 20100 13006 20156
rect 13006 20100 13010 20156
rect 12946 20096 13010 20100
rect 13026 20156 13090 20160
rect 13026 20100 13030 20156
rect 13030 20100 13086 20156
rect 13086 20100 13090 20156
rect 13026 20096 13090 20100
rect 13106 20156 13170 20160
rect 13106 20100 13110 20156
rect 13110 20100 13166 20156
rect 13166 20100 13170 20156
rect 13106 20096 13170 20100
rect 13186 20156 13250 20160
rect 13186 20100 13190 20156
rect 13190 20100 13246 20156
rect 13246 20100 13250 20156
rect 13186 20096 13250 20100
rect 4378 19612 4442 19616
rect 4378 19556 4382 19612
rect 4382 19556 4438 19612
rect 4438 19556 4442 19612
rect 4378 19552 4442 19556
rect 4458 19612 4522 19616
rect 4458 19556 4462 19612
rect 4462 19556 4518 19612
rect 4518 19556 4522 19612
rect 4458 19552 4522 19556
rect 4538 19612 4602 19616
rect 4538 19556 4542 19612
rect 4542 19556 4598 19612
rect 4598 19556 4602 19612
rect 4538 19552 4602 19556
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 7805 19612 7869 19616
rect 7805 19556 7809 19612
rect 7809 19556 7865 19612
rect 7865 19556 7869 19612
rect 7805 19552 7869 19556
rect 7885 19612 7949 19616
rect 7885 19556 7889 19612
rect 7889 19556 7945 19612
rect 7945 19556 7949 19612
rect 7885 19552 7949 19556
rect 7965 19612 8029 19616
rect 7965 19556 7969 19612
rect 7969 19556 8025 19612
rect 8025 19556 8029 19612
rect 7965 19552 8029 19556
rect 8045 19612 8109 19616
rect 8045 19556 8049 19612
rect 8049 19556 8105 19612
rect 8105 19556 8109 19612
rect 8045 19552 8109 19556
rect 11232 19612 11296 19616
rect 11232 19556 11236 19612
rect 11236 19556 11292 19612
rect 11292 19556 11296 19612
rect 11232 19552 11296 19556
rect 11312 19612 11376 19616
rect 11312 19556 11316 19612
rect 11316 19556 11372 19612
rect 11372 19556 11376 19612
rect 11312 19552 11376 19556
rect 11392 19612 11456 19616
rect 11392 19556 11396 19612
rect 11396 19556 11452 19612
rect 11452 19556 11456 19612
rect 11392 19552 11456 19556
rect 11472 19612 11536 19616
rect 11472 19556 11476 19612
rect 11476 19556 11532 19612
rect 11532 19556 11536 19612
rect 11472 19552 11536 19556
rect 14659 19612 14723 19616
rect 14659 19556 14663 19612
rect 14663 19556 14719 19612
rect 14719 19556 14723 19612
rect 14659 19552 14723 19556
rect 14739 19612 14803 19616
rect 14739 19556 14743 19612
rect 14743 19556 14799 19612
rect 14799 19556 14803 19612
rect 14739 19552 14803 19556
rect 14819 19612 14883 19616
rect 14819 19556 14823 19612
rect 14823 19556 14879 19612
rect 14879 19556 14883 19612
rect 14819 19552 14883 19556
rect 14899 19612 14963 19616
rect 14899 19556 14903 19612
rect 14903 19556 14959 19612
rect 14959 19556 14963 19612
rect 14899 19552 14963 19556
rect 2665 19068 2729 19072
rect 2665 19012 2669 19068
rect 2669 19012 2725 19068
rect 2725 19012 2729 19068
rect 2665 19008 2729 19012
rect 2745 19068 2809 19072
rect 2745 19012 2749 19068
rect 2749 19012 2805 19068
rect 2805 19012 2809 19068
rect 2745 19008 2809 19012
rect 2825 19068 2889 19072
rect 2825 19012 2829 19068
rect 2829 19012 2885 19068
rect 2885 19012 2889 19068
rect 2825 19008 2889 19012
rect 2905 19068 2969 19072
rect 2905 19012 2909 19068
rect 2909 19012 2965 19068
rect 2965 19012 2969 19068
rect 2905 19008 2969 19012
rect 6092 19068 6156 19072
rect 6092 19012 6096 19068
rect 6096 19012 6152 19068
rect 6152 19012 6156 19068
rect 6092 19008 6156 19012
rect 6172 19068 6236 19072
rect 6172 19012 6176 19068
rect 6176 19012 6232 19068
rect 6232 19012 6236 19068
rect 6172 19008 6236 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 9519 19068 9583 19072
rect 9519 19012 9523 19068
rect 9523 19012 9579 19068
rect 9579 19012 9583 19068
rect 9519 19008 9583 19012
rect 9599 19068 9663 19072
rect 9599 19012 9603 19068
rect 9603 19012 9659 19068
rect 9659 19012 9663 19068
rect 9599 19008 9663 19012
rect 9679 19068 9743 19072
rect 9679 19012 9683 19068
rect 9683 19012 9739 19068
rect 9739 19012 9743 19068
rect 9679 19008 9743 19012
rect 9759 19068 9823 19072
rect 9759 19012 9763 19068
rect 9763 19012 9819 19068
rect 9819 19012 9823 19068
rect 9759 19008 9823 19012
rect 12946 19068 13010 19072
rect 12946 19012 12950 19068
rect 12950 19012 13006 19068
rect 13006 19012 13010 19068
rect 12946 19008 13010 19012
rect 13026 19068 13090 19072
rect 13026 19012 13030 19068
rect 13030 19012 13086 19068
rect 13086 19012 13090 19068
rect 13026 19008 13090 19012
rect 13106 19068 13170 19072
rect 13106 19012 13110 19068
rect 13110 19012 13166 19068
rect 13166 19012 13170 19068
rect 13106 19008 13170 19012
rect 13186 19068 13250 19072
rect 13186 19012 13190 19068
rect 13190 19012 13246 19068
rect 13246 19012 13250 19068
rect 13186 19008 13250 19012
rect 4378 18524 4442 18528
rect 4378 18468 4382 18524
rect 4382 18468 4438 18524
rect 4438 18468 4442 18524
rect 4378 18464 4442 18468
rect 4458 18524 4522 18528
rect 4458 18468 4462 18524
rect 4462 18468 4518 18524
rect 4518 18468 4522 18524
rect 4458 18464 4522 18468
rect 4538 18524 4602 18528
rect 4538 18468 4542 18524
rect 4542 18468 4598 18524
rect 4598 18468 4602 18524
rect 4538 18464 4602 18468
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 7805 18524 7869 18528
rect 7805 18468 7809 18524
rect 7809 18468 7865 18524
rect 7865 18468 7869 18524
rect 7805 18464 7869 18468
rect 7885 18524 7949 18528
rect 7885 18468 7889 18524
rect 7889 18468 7945 18524
rect 7945 18468 7949 18524
rect 7885 18464 7949 18468
rect 7965 18524 8029 18528
rect 7965 18468 7969 18524
rect 7969 18468 8025 18524
rect 8025 18468 8029 18524
rect 7965 18464 8029 18468
rect 8045 18524 8109 18528
rect 8045 18468 8049 18524
rect 8049 18468 8105 18524
rect 8105 18468 8109 18524
rect 8045 18464 8109 18468
rect 11232 18524 11296 18528
rect 11232 18468 11236 18524
rect 11236 18468 11292 18524
rect 11292 18468 11296 18524
rect 11232 18464 11296 18468
rect 11312 18524 11376 18528
rect 11312 18468 11316 18524
rect 11316 18468 11372 18524
rect 11372 18468 11376 18524
rect 11312 18464 11376 18468
rect 11392 18524 11456 18528
rect 11392 18468 11396 18524
rect 11396 18468 11452 18524
rect 11452 18468 11456 18524
rect 11392 18464 11456 18468
rect 11472 18524 11536 18528
rect 11472 18468 11476 18524
rect 11476 18468 11532 18524
rect 11532 18468 11536 18524
rect 11472 18464 11536 18468
rect 14659 18524 14723 18528
rect 14659 18468 14663 18524
rect 14663 18468 14719 18524
rect 14719 18468 14723 18524
rect 14659 18464 14723 18468
rect 14739 18524 14803 18528
rect 14739 18468 14743 18524
rect 14743 18468 14799 18524
rect 14799 18468 14803 18524
rect 14739 18464 14803 18468
rect 14819 18524 14883 18528
rect 14819 18468 14823 18524
rect 14823 18468 14879 18524
rect 14879 18468 14883 18524
rect 14819 18464 14883 18468
rect 14899 18524 14963 18528
rect 14899 18468 14903 18524
rect 14903 18468 14959 18524
rect 14959 18468 14963 18524
rect 14899 18464 14963 18468
rect 2665 17980 2729 17984
rect 2665 17924 2669 17980
rect 2669 17924 2725 17980
rect 2725 17924 2729 17980
rect 2665 17920 2729 17924
rect 2745 17980 2809 17984
rect 2745 17924 2749 17980
rect 2749 17924 2805 17980
rect 2805 17924 2809 17980
rect 2745 17920 2809 17924
rect 2825 17980 2889 17984
rect 2825 17924 2829 17980
rect 2829 17924 2885 17980
rect 2885 17924 2889 17980
rect 2825 17920 2889 17924
rect 2905 17980 2969 17984
rect 2905 17924 2909 17980
rect 2909 17924 2965 17980
rect 2965 17924 2969 17980
rect 2905 17920 2969 17924
rect 6092 17980 6156 17984
rect 6092 17924 6096 17980
rect 6096 17924 6152 17980
rect 6152 17924 6156 17980
rect 6092 17920 6156 17924
rect 6172 17980 6236 17984
rect 6172 17924 6176 17980
rect 6176 17924 6232 17980
rect 6232 17924 6236 17980
rect 6172 17920 6236 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 9519 17980 9583 17984
rect 9519 17924 9523 17980
rect 9523 17924 9579 17980
rect 9579 17924 9583 17980
rect 9519 17920 9583 17924
rect 9599 17980 9663 17984
rect 9599 17924 9603 17980
rect 9603 17924 9659 17980
rect 9659 17924 9663 17980
rect 9599 17920 9663 17924
rect 9679 17980 9743 17984
rect 9679 17924 9683 17980
rect 9683 17924 9739 17980
rect 9739 17924 9743 17980
rect 9679 17920 9743 17924
rect 9759 17980 9823 17984
rect 9759 17924 9763 17980
rect 9763 17924 9819 17980
rect 9819 17924 9823 17980
rect 9759 17920 9823 17924
rect 12946 17980 13010 17984
rect 12946 17924 12950 17980
rect 12950 17924 13006 17980
rect 13006 17924 13010 17980
rect 12946 17920 13010 17924
rect 13026 17980 13090 17984
rect 13026 17924 13030 17980
rect 13030 17924 13086 17980
rect 13086 17924 13090 17980
rect 13026 17920 13090 17924
rect 13106 17980 13170 17984
rect 13106 17924 13110 17980
rect 13110 17924 13166 17980
rect 13166 17924 13170 17980
rect 13106 17920 13170 17924
rect 13186 17980 13250 17984
rect 13186 17924 13190 17980
rect 13190 17924 13246 17980
rect 13246 17924 13250 17980
rect 13186 17920 13250 17924
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 45184 2977 45744
rect 2657 45120 2665 45184
rect 2729 45120 2745 45184
rect 2809 45120 2825 45184
rect 2889 45120 2905 45184
rect 2969 45120 2977 45184
rect 2657 44096 2977 45120
rect 2657 44032 2665 44096
rect 2729 44032 2745 44096
rect 2809 44032 2825 44096
rect 2889 44032 2905 44096
rect 2969 44032 2977 44096
rect 2657 43008 2977 44032
rect 2657 42944 2665 43008
rect 2729 42944 2745 43008
rect 2809 42944 2825 43008
rect 2889 42944 2905 43008
rect 2969 42944 2977 43008
rect 2657 41920 2977 42944
rect 2657 41856 2665 41920
rect 2729 41856 2745 41920
rect 2809 41856 2825 41920
rect 2889 41856 2905 41920
rect 2969 41856 2977 41920
rect 2657 40832 2977 41856
rect 2657 40768 2665 40832
rect 2729 40768 2745 40832
rect 2809 40768 2825 40832
rect 2889 40768 2905 40832
rect 2969 40768 2977 40832
rect 2657 39744 2977 40768
rect 2657 39680 2665 39744
rect 2729 39680 2745 39744
rect 2809 39680 2825 39744
rect 2889 39680 2905 39744
rect 2969 39680 2977 39744
rect 2657 38656 2977 39680
rect 2657 38592 2665 38656
rect 2729 38592 2745 38656
rect 2809 38592 2825 38656
rect 2889 38592 2905 38656
rect 2969 38592 2977 38656
rect 2657 37568 2977 38592
rect 2657 37504 2665 37568
rect 2729 37504 2745 37568
rect 2809 37504 2825 37568
rect 2889 37504 2905 37568
rect 2969 37504 2977 37568
rect 2657 36480 2977 37504
rect 2657 36416 2665 36480
rect 2729 36416 2745 36480
rect 2809 36416 2825 36480
rect 2889 36416 2905 36480
rect 2969 36416 2977 36480
rect 2657 35392 2977 36416
rect 2657 35328 2665 35392
rect 2729 35328 2745 35392
rect 2809 35328 2825 35392
rect 2889 35328 2905 35392
rect 2969 35328 2977 35392
rect 2657 34304 2977 35328
rect 2657 34240 2665 34304
rect 2729 34240 2745 34304
rect 2809 34240 2825 34304
rect 2889 34240 2905 34304
rect 2969 34240 2977 34304
rect 2657 33216 2977 34240
rect 2657 33152 2665 33216
rect 2729 33152 2745 33216
rect 2809 33152 2825 33216
rect 2889 33152 2905 33216
rect 2969 33152 2977 33216
rect 2657 32128 2977 33152
rect 2657 32064 2665 32128
rect 2729 32064 2745 32128
rect 2809 32064 2825 32128
rect 2889 32064 2905 32128
rect 2969 32064 2977 32128
rect 2657 31040 2977 32064
rect 2657 30976 2665 31040
rect 2729 30976 2745 31040
rect 2809 30976 2825 31040
rect 2889 30976 2905 31040
rect 2969 30976 2977 31040
rect 2657 29952 2977 30976
rect 2657 29888 2665 29952
rect 2729 29888 2745 29952
rect 2809 29888 2825 29952
rect 2889 29888 2905 29952
rect 2969 29888 2977 29952
rect 2657 28864 2977 29888
rect 2657 28800 2665 28864
rect 2729 28800 2745 28864
rect 2809 28800 2825 28864
rect 2889 28800 2905 28864
rect 2969 28800 2977 28864
rect 2657 27776 2977 28800
rect 2657 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2977 27776
rect 2657 26688 2977 27712
rect 2657 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2977 26688
rect 2657 25600 2977 26624
rect 2657 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2977 25600
rect 2657 24512 2977 25536
rect 2657 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2977 24512
rect 2657 23424 2977 24448
rect 2657 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2977 23424
rect 2657 22336 2977 23360
rect 2657 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2977 22336
rect 2657 21248 2977 22272
rect 2657 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2977 21248
rect 2657 20160 2977 21184
rect 2657 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2977 20160
rect 2657 19072 2977 20096
rect 2657 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2977 19072
rect 2657 17984 2977 19008
rect 2657 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2977 17984
rect 2657 16896 2977 17920
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 45728 4690 45744
rect 4370 45664 4378 45728
rect 4442 45664 4458 45728
rect 4522 45664 4538 45728
rect 4602 45664 4618 45728
rect 4682 45664 4690 45728
rect 4370 44640 4690 45664
rect 4370 44576 4378 44640
rect 4442 44576 4458 44640
rect 4522 44576 4538 44640
rect 4602 44576 4618 44640
rect 4682 44576 4690 44640
rect 4370 43552 4690 44576
rect 4370 43488 4378 43552
rect 4442 43488 4458 43552
rect 4522 43488 4538 43552
rect 4602 43488 4618 43552
rect 4682 43488 4690 43552
rect 4370 42464 4690 43488
rect 4370 42400 4378 42464
rect 4442 42400 4458 42464
rect 4522 42400 4538 42464
rect 4602 42400 4618 42464
rect 4682 42400 4690 42464
rect 4370 41376 4690 42400
rect 4370 41312 4378 41376
rect 4442 41312 4458 41376
rect 4522 41312 4538 41376
rect 4602 41312 4618 41376
rect 4682 41312 4690 41376
rect 4370 40288 4690 41312
rect 4370 40224 4378 40288
rect 4442 40224 4458 40288
rect 4522 40224 4538 40288
rect 4602 40224 4618 40288
rect 4682 40224 4690 40288
rect 4370 39200 4690 40224
rect 4370 39136 4378 39200
rect 4442 39136 4458 39200
rect 4522 39136 4538 39200
rect 4602 39136 4618 39200
rect 4682 39136 4690 39200
rect 4370 38112 4690 39136
rect 4370 38048 4378 38112
rect 4442 38048 4458 38112
rect 4522 38048 4538 38112
rect 4602 38048 4618 38112
rect 4682 38048 4690 38112
rect 4370 37024 4690 38048
rect 4370 36960 4378 37024
rect 4442 36960 4458 37024
rect 4522 36960 4538 37024
rect 4602 36960 4618 37024
rect 4682 36960 4690 37024
rect 4370 35936 4690 36960
rect 4370 35872 4378 35936
rect 4442 35872 4458 35936
rect 4522 35872 4538 35936
rect 4602 35872 4618 35936
rect 4682 35872 4690 35936
rect 4370 34848 4690 35872
rect 4370 34784 4378 34848
rect 4442 34784 4458 34848
rect 4522 34784 4538 34848
rect 4602 34784 4618 34848
rect 4682 34784 4690 34848
rect 4370 33760 4690 34784
rect 4370 33696 4378 33760
rect 4442 33696 4458 33760
rect 4522 33696 4538 33760
rect 4602 33696 4618 33760
rect 4682 33696 4690 33760
rect 4370 32672 4690 33696
rect 4370 32608 4378 32672
rect 4442 32608 4458 32672
rect 4522 32608 4538 32672
rect 4602 32608 4618 32672
rect 4682 32608 4690 32672
rect 4370 31584 4690 32608
rect 4370 31520 4378 31584
rect 4442 31520 4458 31584
rect 4522 31520 4538 31584
rect 4602 31520 4618 31584
rect 4682 31520 4690 31584
rect 4370 30496 4690 31520
rect 4370 30432 4378 30496
rect 4442 30432 4458 30496
rect 4522 30432 4538 30496
rect 4602 30432 4618 30496
rect 4682 30432 4690 30496
rect 4370 29408 4690 30432
rect 4370 29344 4378 29408
rect 4442 29344 4458 29408
rect 4522 29344 4538 29408
rect 4602 29344 4618 29408
rect 4682 29344 4690 29408
rect 4370 28320 4690 29344
rect 4370 28256 4378 28320
rect 4442 28256 4458 28320
rect 4522 28256 4538 28320
rect 4602 28256 4618 28320
rect 4682 28256 4690 28320
rect 4370 27232 4690 28256
rect 4370 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4690 27232
rect 4370 26144 4690 27168
rect 4370 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4690 26144
rect 4370 25056 4690 26080
rect 4370 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4690 25056
rect 4370 23968 4690 24992
rect 4370 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4690 23968
rect 4370 22880 4690 23904
rect 4370 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4690 22880
rect 4370 21792 4690 22816
rect 4370 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4690 21792
rect 4370 20704 4690 21728
rect 4370 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4690 20704
rect 4370 19616 4690 20640
rect 4370 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4690 19616
rect 4370 18528 4690 19552
rect 4370 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4690 18528
rect 4370 17440 4690 18464
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 45184 6404 45744
rect 6084 45120 6092 45184
rect 6156 45120 6172 45184
rect 6236 45120 6252 45184
rect 6316 45120 6332 45184
rect 6396 45120 6404 45184
rect 6084 44096 6404 45120
rect 6084 44032 6092 44096
rect 6156 44032 6172 44096
rect 6236 44032 6252 44096
rect 6316 44032 6332 44096
rect 6396 44032 6404 44096
rect 6084 43008 6404 44032
rect 6084 42944 6092 43008
rect 6156 42944 6172 43008
rect 6236 42944 6252 43008
rect 6316 42944 6332 43008
rect 6396 42944 6404 43008
rect 6084 41920 6404 42944
rect 6084 41856 6092 41920
rect 6156 41856 6172 41920
rect 6236 41856 6252 41920
rect 6316 41856 6332 41920
rect 6396 41856 6404 41920
rect 6084 40832 6404 41856
rect 6084 40768 6092 40832
rect 6156 40768 6172 40832
rect 6236 40768 6252 40832
rect 6316 40768 6332 40832
rect 6396 40768 6404 40832
rect 6084 39744 6404 40768
rect 6084 39680 6092 39744
rect 6156 39680 6172 39744
rect 6236 39680 6252 39744
rect 6316 39680 6332 39744
rect 6396 39680 6404 39744
rect 6084 38656 6404 39680
rect 6084 38592 6092 38656
rect 6156 38592 6172 38656
rect 6236 38592 6252 38656
rect 6316 38592 6332 38656
rect 6396 38592 6404 38656
rect 6084 37568 6404 38592
rect 6084 37504 6092 37568
rect 6156 37504 6172 37568
rect 6236 37504 6252 37568
rect 6316 37504 6332 37568
rect 6396 37504 6404 37568
rect 6084 36480 6404 37504
rect 6084 36416 6092 36480
rect 6156 36416 6172 36480
rect 6236 36416 6252 36480
rect 6316 36416 6332 36480
rect 6396 36416 6404 36480
rect 6084 35392 6404 36416
rect 6084 35328 6092 35392
rect 6156 35328 6172 35392
rect 6236 35328 6252 35392
rect 6316 35328 6332 35392
rect 6396 35328 6404 35392
rect 6084 34304 6404 35328
rect 6084 34240 6092 34304
rect 6156 34240 6172 34304
rect 6236 34240 6252 34304
rect 6316 34240 6332 34304
rect 6396 34240 6404 34304
rect 6084 33216 6404 34240
rect 6084 33152 6092 33216
rect 6156 33152 6172 33216
rect 6236 33152 6252 33216
rect 6316 33152 6332 33216
rect 6396 33152 6404 33216
rect 6084 32128 6404 33152
rect 6084 32064 6092 32128
rect 6156 32064 6172 32128
rect 6236 32064 6252 32128
rect 6316 32064 6332 32128
rect 6396 32064 6404 32128
rect 6084 31040 6404 32064
rect 6084 30976 6092 31040
rect 6156 30976 6172 31040
rect 6236 30976 6252 31040
rect 6316 30976 6332 31040
rect 6396 30976 6404 31040
rect 6084 29952 6404 30976
rect 6084 29888 6092 29952
rect 6156 29888 6172 29952
rect 6236 29888 6252 29952
rect 6316 29888 6332 29952
rect 6396 29888 6404 29952
rect 6084 28864 6404 29888
rect 6084 28800 6092 28864
rect 6156 28800 6172 28864
rect 6236 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6404 28864
rect 6084 27776 6404 28800
rect 6084 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6404 27776
rect 6084 26688 6404 27712
rect 6084 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6404 26688
rect 6084 25600 6404 26624
rect 6084 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6404 25600
rect 6084 24512 6404 25536
rect 6084 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6404 24512
rect 6084 23424 6404 24448
rect 6084 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6404 23424
rect 6084 22336 6404 23360
rect 6084 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6404 22336
rect 6084 21248 6404 22272
rect 6084 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6404 21248
rect 6084 20160 6404 21184
rect 6084 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6404 20160
rect 6084 19072 6404 20096
rect 6084 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6404 19072
rect 6084 17984 6404 19008
rect 6084 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6404 17984
rect 6084 16896 6404 17920
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 45728 8117 45744
rect 7797 45664 7805 45728
rect 7869 45664 7885 45728
rect 7949 45664 7965 45728
rect 8029 45664 8045 45728
rect 8109 45664 8117 45728
rect 7797 44640 8117 45664
rect 7797 44576 7805 44640
rect 7869 44576 7885 44640
rect 7949 44576 7965 44640
rect 8029 44576 8045 44640
rect 8109 44576 8117 44640
rect 7797 43552 8117 44576
rect 7797 43488 7805 43552
rect 7869 43488 7885 43552
rect 7949 43488 7965 43552
rect 8029 43488 8045 43552
rect 8109 43488 8117 43552
rect 7797 42464 8117 43488
rect 7797 42400 7805 42464
rect 7869 42400 7885 42464
rect 7949 42400 7965 42464
rect 8029 42400 8045 42464
rect 8109 42400 8117 42464
rect 7797 41376 8117 42400
rect 7797 41312 7805 41376
rect 7869 41312 7885 41376
rect 7949 41312 7965 41376
rect 8029 41312 8045 41376
rect 8109 41312 8117 41376
rect 7797 40288 8117 41312
rect 7797 40224 7805 40288
rect 7869 40224 7885 40288
rect 7949 40224 7965 40288
rect 8029 40224 8045 40288
rect 8109 40224 8117 40288
rect 7797 39200 8117 40224
rect 7797 39136 7805 39200
rect 7869 39136 7885 39200
rect 7949 39136 7965 39200
rect 8029 39136 8045 39200
rect 8109 39136 8117 39200
rect 7797 38112 8117 39136
rect 7797 38048 7805 38112
rect 7869 38048 7885 38112
rect 7949 38048 7965 38112
rect 8029 38048 8045 38112
rect 8109 38048 8117 38112
rect 7797 37024 8117 38048
rect 7797 36960 7805 37024
rect 7869 36960 7885 37024
rect 7949 36960 7965 37024
rect 8029 36960 8045 37024
rect 8109 36960 8117 37024
rect 7797 35936 8117 36960
rect 7797 35872 7805 35936
rect 7869 35872 7885 35936
rect 7949 35872 7965 35936
rect 8029 35872 8045 35936
rect 8109 35872 8117 35936
rect 7797 34848 8117 35872
rect 7797 34784 7805 34848
rect 7869 34784 7885 34848
rect 7949 34784 7965 34848
rect 8029 34784 8045 34848
rect 8109 34784 8117 34848
rect 7797 33760 8117 34784
rect 7797 33696 7805 33760
rect 7869 33696 7885 33760
rect 7949 33696 7965 33760
rect 8029 33696 8045 33760
rect 8109 33696 8117 33760
rect 7797 32672 8117 33696
rect 7797 32608 7805 32672
rect 7869 32608 7885 32672
rect 7949 32608 7965 32672
rect 8029 32608 8045 32672
rect 8109 32608 8117 32672
rect 7797 31584 8117 32608
rect 7797 31520 7805 31584
rect 7869 31520 7885 31584
rect 7949 31520 7965 31584
rect 8029 31520 8045 31584
rect 8109 31520 8117 31584
rect 7797 30496 8117 31520
rect 7797 30432 7805 30496
rect 7869 30432 7885 30496
rect 7949 30432 7965 30496
rect 8029 30432 8045 30496
rect 8109 30432 8117 30496
rect 7797 29408 8117 30432
rect 7797 29344 7805 29408
rect 7869 29344 7885 29408
rect 7949 29344 7965 29408
rect 8029 29344 8045 29408
rect 8109 29344 8117 29408
rect 7797 28320 8117 29344
rect 7797 28256 7805 28320
rect 7869 28256 7885 28320
rect 7949 28256 7965 28320
rect 8029 28256 8045 28320
rect 8109 28256 8117 28320
rect 7797 27232 8117 28256
rect 7797 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8117 27232
rect 7797 26144 8117 27168
rect 7797 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8117 26144
rect 7797 25056 8117 26080
rect 7797 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8117 25056
rect 7797 23968 8117 24992
rect 7797 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8117 23968
rect 7797 22880 8117 23904
rect 7797 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8117 22880
rect 7797 21792 8117 22816
rect 7797 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8117 21792
rect 7797 20704 8117 21728
rect 7797 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8117 20704
rect 7797 19616 8117 20640
rect 7797 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8117 19616
rect 7797 18528 8117 19552
rect 7797 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8117 18528
rect 7797 17440 8117 18464
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 45184 9831 45744
rect 9511 45120 9519 45184
rect 9583 45120 9599 45184
rect 9663 45120 9679 45184
rect 9743 45120 9759 45184
rect 9823 45120 9831 45184
rect 9511 44096 9831 45120
rect 9511 44032 9519 44096
rect 9583 44032 9599 44096
rect 9663 44032 9679 44096
rect 9743 44032 9759 44096
rect 9823 44032 9831 44096
rect 9511 43008 9831 44032
rect 9511 42944 9519 43008
rect 9583 42944 9599 43008
rect 9663 42944 9679 43008
rect 9743 42944 9759 43008
rect 9823 42944 9831 43008
rect 9511 41920 9831 42944
rect 9511 41856 9519 41920
rect 9583 41856 9599 41920
rect 9663 41856 9679 41920
rect 9743 41856 9759 41920
rect 9823 41856 9831 41920
rect 9511 40832 9831 41856
rect 9511 40768 9519 40832
rect 9583 40768 9599 40832
rect 9663 40768 9679 40832
rect 9743 40768 9759 40832
rect 9823 40768 9831 40832
rect 9511 39744 9831 40768
rect 9511 39680 9519 39744
rect 9583 39680 9599 39744
rect 9663 39680 9679 39744
rect 9743 39680 9759 39744
rect 9823 39680 9831 39744
rect 9511 38656 9831 39680
rect 9511 38592 9519 38656
rect 9583 38592 9599 38656
rect 9663 38592 9679 38656
rect 9743 38592 9759 38656
rect 9823 38592 9831 38656
rect 9511 37568 9831 38592
rect 9511 37504 9519 37568
rect 9583 37504 9599 37568
rect 9663 37504 9679 37568
rect 9743 37504 9759 37568
rect 9823 37504 9831 37568
rect 9511 36480 9831 37504
rect 9511 36416 9519 36480
rect 9583 36416 9599 36480
rect 9663 36416 9679 36480
rect 9743 36416 9759 36480
rect 9823 36416 9831 36480
rect 9511 35392 9831 36416
rect 9511 35328 9519 35392
rect 9583 35328 9599 35392
rect 9663 35328 9679 35392
rect 9743 35328 9759 35392
rect 9823 35328 9831 35392
rect 9511 34304 9831 35328
rect 9511 34240 9519 34304
rect 9583 34240 9599 34304
rect 9663 34240 9679 34304
rect 9743 34240 9759 34304
rect 9823 34240 9831 34304
rect 9511 33216 9831 34240
rect 9511 33152 9519 33216
rect 9583 33152 9599 33216
rect 9663 33152 9679 33216
rect 9743 33152 9759 33216
rect 9823 33152 9831 33216
rect 9511 32128 9831 33152
rect 9511 32064 9519 32128
rect 9583 32064 9599 32128
rect 9663 32064 9679 32128
rect 9743 32064 9759 32128
rect 9823 32064 9831 32128
rect 9511 31040 9831 32064
rect 9511 30976 9519 31040
rect 9583 30976 9599 31040
rect 9663 30976 9679 31040
rect 9743 30976 9759 31040
rect 9823 30976 9831 31040
rect 9511 29952 9831 30976
rect 9511 29888 9519 29952
rect 9583 29888 9599 29952
rect 9663 29888 9679 29952
rect 9743 29888 9759 29952
rect 9823 29888 9831 29952
rect 9511 28864 9831 29888
rect 9511 28800 9519 28864
rect 9583 28800 9599 28864
rect 9663 28800 9679 28864
rect 9743 28800 9759 28864
rect 9823 28800 9831 28864
rect 9511 27776 9831 28800
rect 9511 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9831 27776
rect 9511 26688 9831 27712
rect 9511 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9831 26688
rect 9511 25600 9831 26624
rect 9511 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9831 25600
rect 9511 24512 9831 25536
rect 9511 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9831 24512
rect 9511 23424 9831 24448
rect 9511 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9831 23424
rect 9511 22336 9831 23360
rect 9511 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9831 22336
rect 9511 21248 9831 22272
rect 9511 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9831 21248
rect 9511 20160 9831 21184
rect 9511 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9831 20160
rect 9511 19072 9831 20096
rect 9511 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9831 19072
rect 9511 17984 9831 19008
rect 9511 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9831 17984
rect 9511 16896 9831 17920
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 45728 11544 45744
rect 11224 45664 11232 45728
rect 11296 45664 11312 45728
rect 11376 45664 11392 45728
rect 11456 45664 11472 45728
rect 11536 45664 11544 45728
rect 11224 44640 11544 45664
rect 11224 44576 11232 44640
rect 11296 44576 11312 44640
rect 11376 44576 11392 44640
rect 11456 44576 11472 44640
rect 11536 44576 11544 44640
rect 11224 43552 11544 44576
rect 11224 43488 11232 43552
rect 11296 43488 11312 43552
rect 11376 43488 11392 43552
rect 11456 43488 11472 43552
rect 11536 43488 11544 43552
rect 11224 42464 11544 43488
rect 11224 42400 11232 42464
rect 11296 42400 11312 42464
rect 11376 42400 11392 42464
rect 11456 42400 11472 42464
rect 11536 42400 11544 42464
rect 11224 41376 11544 42400
rect 11224 41312 11232 41376
rect 11296 41312 11312 41376
rect 11376 41312 11392 41376
rect 11456 41312 11472 41376
rect 11536 41312 11544 41376
rect 11224 40288 11544 41312
rect 11224 40224 11232 40288
rect 11296 40224 11312 40288
rect 11376 40224 11392 40288
rect 11456 40224 11472 40288
rect 11536 40224 11544 40288
rect 11224 39200 11544 40224
rect 11224 39136 11232 39200
rect 11296 39136 11312 39200
rect 11376 39136 11392 39200
rect 11456 39136 11472 39200
rect 11536 39136 11544 39200
rect 11224 38112 11544 39136
rect 11224 38048 11232 38112
rect 11296 38048 11312 38112
rect 11376 38048 11392 38112
rect 11456 38048 11472 38112
rect 11536 38048 11544 38112
rect 11224 37024 11544 38048
rect 11224 36960 11232 37024
rect 11296 36960 11312 37024
rect 11376 36960 11392 37024
rect 11456 36960 11472 37024
rect 11536 36960 11544 37024
rect 11224 35936 11544 36960
rect 11224 35872 11232 35936
rect 11296 35872 11312 35936
rect 11376 35872 11392 35936
rect 11456 35872 11472 35936
rect 11536 35872 11544 35936
rect 11224 34848 11544 35872
rect 11224 34784 11232 34848
rect 11296 34784 11312 34848
rect 11376 34784 11392 34848
rect 11456 34784 11472 34848
rect 11536 34784 11544 34848
rect 11224 33760 11544 34784
rect 11224 33696 11232 33760
rect 11296 33696 11312 33760
rect 11376 33696 11392 33760
rect 11456 33696 11472 33760
rect 11536 33696 11544 33760
rect 11224 32672 11544 33696
rect 11224 32608 11232 32672
rect 11296 32608 11312 32672
rect 11376 32608 11392 32672
rect 11456 32608 11472 32672
rect 11536 32608 11544 32672
rect 11224 31584 11544 32608
rect 11224 31520 11232 31584
rect 11296 31520 11312 31584
rect 11376 31520 11392 31584
rect 11456 31520 11472 31584
rect 11536 31520 11544 31584
rect 11224 30496 11544 31520
rect 11224 30432 11232 30496
rect 11296 30432 11312 30496
rect 11376 30432 11392 30496
rect 11456 30432 11472 30496
rect 11536 30432 11544 30496
rect 11224 29408 11544 30432
rect 11224 29344 11232 29408
rect 11296 29344 11312 29408
rect 11376 29344 11392 29408
rect 11456 29344 11472 29408
rect 11536 29344 11544 29408
rect 11224 28320 11544 29344
rect 11224 28256 11232 28320
rect 11296 28256 11312 28320
rect 11376 28256 11392 28320
rect 11456 28256 11472 28320
rect 11536 28256 11544 28320
rect 11224 27232 11544 28256
rect 11224 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11544 27232
rect 11224 26144 11544 27168
rect 11224 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11544 26144
rect 11224 25056 11544 26080
rect 11224 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11544 25056
rect 11224 23968 11544 24992
rect 11224 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11544 23968
rect 11224 22880 11544 23904
rect 11224 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11544 22880
rect 11224 21792 11544 22816
rect 11224 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11544 21792
rect 11224 20704 11544 21728
rect 11224 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11544 20704
rect 11224 19616 11544 20640
rect 11224 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11544 19616
rect 11224 18528 11544 19552
rect 11224 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11544 18528
rect 11224 17440 11544 18464
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 45184 13258 45744
rect 12938 45120 12946 45184
rect 13010 45120 13026 45184
rect 13090 45120 13106 45184
rect 13170 45120 13186 45184
rect 13250 45120 13258 45184
rect 12938 44096 13258 45120
rect 12938 44032 12946 44096
rect 13010 44032 13026 44096
rect 13090 44032 13106 44096
rect 13170 44032 13186 44096
rect 13250 44032 13258 44096
rect 12938 43008 13258 44032
rect 12938 42944 12946 43008
rect 13010 42944 13026 43008
rect 13090 42944 13106 43008
rect 13170 42944 13186 43008
rect 13250 42944 13258 43008
rect 12938 41920 13258 42944
rect 12938 41856 12946 41920
rect 13010 41856 13026 41920
rect 13090 41856 13106 41920
rect 13170 41856 13186 41920
rect 13250 41856 13258 41920
rect 12938 40832 13258 41856
rect 12938 40768 12946 40832
rect 13010 40768 13026 40832
rect 13090 40768 13106 40832
rect 13170 40768 13186 40832
rect 13250 40768 13258 40832
rect 12938 39744 13258 40768
rect 12938 39680 12946 39744
rect 13010 39680 13026 39744
rect 13090 39680 13106 39744
rect 13170 39680 13186 39744
rect 13250 39680 13258 39744
rect 12938 38656 13258 39680
rect 12938 38592 12946 38656
rect 13010 38592 13026 38656
rect 13090 38592 13106 38656
rect 13170 38592 13186 38656
rect 13250 38592 13258 38656
rect 12938 37568 13258 38592
rect 12938 37504 12946 37568
rect 13010 37504 13026 37568
rect 13090 37504 13106 37568
rect 13170 37504 13186 37568
rect 13250 37504 13258 37568
rect 12938 36480 13258 37504
rect 12938 36416 12946 36480
rect 13010 36416 13026 36480
rect 13090 36416 13106 36480
rect 13170 36416 13186 36480
rect 13250 36416 13258 36480
rect 12938 35392 13258 36416
rect 12938 35328 12946 35392
rect 13010 35328 13026 35392
rect 13090 35328 13106 35392
rect 13170 35328 13186 35392
rect 13250 35328 13258 35392
rect 12938 34304 13258 35328
rect 12938 34240 12946 34304
rect 13010 34240 13026 34304
rect 13090 34240 13106 34304
rect 13170 34240 13186 34304
rect 13250 34240 13258 34304
rect 12938 33216 13258 34240
rect 12938 33152 12946 33216
rect 13010 33152 13026 33216
rect 13090 33152 13106 33216
rect 13170 33152 13186 33216
rect 13250 33152 13258 33216
rect 12938 32128 13258 33152
rect 12938 32064 12946 32128
rect 13010 32064 13026 32128
rect 13090 32064 13106 32128
rect 13170 32064 13186 32128
rect 13250 32064 13258 32128
rect 12938 31040 13258 32064
rect 12938 30976 12946 31040
rect 13010 30976 13026 31040
rect 13090 30976 13106 31040
rect 13170 30976 13186 31040
rect 13250 30976 13258 31040
rect 12938 29952 13258 30976
rect 12938 29888 12946 29952
rect 13010 29888 13026 29952
rect 13090 29888 13106 29952
rect 13170 29888 13186 29952
rect 13250 29888 13258 29952
rect 12938 28864 13258 29888
rect 12938 28800 12946 28864
rect 13010 28800 13026 28864
rect 13090 28800 13106 28864
rect 13170 28800 13186 28864
rect 13250 28800 13258 28864
rect 12938 27776 13258 28800
rect 12938 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13258 27776
rect 12938 26688 13258 27712
rect 12938 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13258 26688
rect 12938 25600 13258 26624
rect 12938 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13258 25600
rect 12938 24512 13258 25536
rect 12938 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13258 24512
rect 12938 23424 13258 24448
rect 12938 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13258 23424
rect 12938 22336 13258 23360
rect 12938 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13258 22336
rect 12938 21248 13258 22272
rect 12938 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13258 21248
rect 12938 20160 13258 21184
rect 12938 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13258 20160
rect 12938 19072 13258 20096
rect 12938 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13258 19072
rect 12938 17984 13258 19008
rect 12938 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13258 17984
rect 12938 16896 13258 17920
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 45728 14971 45744
rect 14651 45664 14659 45728
rect 14723 45664 14739 45728
rect 14803 45664 14819 45728
rect 14883 45664 14899 45728
rect 14963 45664 14971 45728
rect 14651 44640 14971 45664
rect 14651 44576 14659 44640
rect 14723 44576 14739 44640
rect 14803 44576 14819 44640
rect 14883 44576 14899 44640
rect 14963 44576 14971 44640
rect 14651 43552 14971 44576
rect 14651 43488 14659 43552
rect 14723 43488 14739 43552
rect 14803 43488 14819 43552
rect 14883 43488 14899 43552
rect 14963 43488 14971 43552
rect 14651 42464 14971 43488
rect 14651 42400 14659 42464
rect 14723 42400 14739 42464
rect 14803 42400 14819 42464
rect 14883 42400 14899 42464
rect 14963 42400 14971 42464
rect 14651 41376 14971 42400
rect 14651 41312 14659 41376
rect 14723 41312 14739 41376
rect 14803 41312 14819 41376
rect 14883 41312 14899 41376
rect 14963 41312 14971 41376
rect 14651 40288 14971 41312
rect 14651 40224 14659 40288
rect 14723 40224 14739 40288
rect 14803 40224 14819 40288
rect 14883 40224 14899 40288
rect 14963 40224 14971 40288
rect 14651 39200 14971 40224
rect 14651 39136 14659 39200
rect 14723 39136 14739 39200
rect 14803 39136 14819 39200
rect 14883 39136 14899 39200
rect 14963 39136 14971 39200
rect 14651 38112 14971 39136
rect 14651 38048 14659 38112
rect 14723 38048 14739 38112
rect 14803 38048 14819 38112
rect 14883 38048 14899 38112
rect 14963 38048 14971 38112
rect 14651 37024 14971 38048
rect 14651 36960 14659 37024
rect 14723 36960 14739 37024
rect 14803 36960 14819 37024
rect 14883 36960 14899 37024
rect 14963 36960 14971 37024
rect 14651 35936 14971 36960
rect 14651 35872 14659 35936
rect 14723 35872 14739 35936
rect 14803 35872 14819 35936
rect 14883 35872 14899 35936
rect 14963 35872 14971 35936
rect 14651 34848 14971 35872
rect 14651 34784 14659 34848
rect 14723 34784 14739 34848
rect 14803 34784 14819 34848
rect 14883 34784 14899 34848
rect 14963 34784 14971 34848
rect 14651 33760 14971 34784
rect 14651 33696 14659 33760
rect 14723 33696 14739 33760
rect 14803 33696 14819 33760
rect 14883 33696 14899 33760
rect 14963 33696 14971 33760
rect 14651 32672 14971 33696
rect 14651 32608 14659 32672
rect 14723 32608 14739 32672
rect 14803 32608 14819 32672
rect 14883 32608 14899 32672
rect 14963 32608 14971 32672
rect 14651 31584 14971 32608
rect 14651 31520 14659 31584
rect 14723 31520 14739 31584
rect 14803 31520 14819 31584
rect 14883 31520 14899 31584
rect 14963 31520 14971 31584
rect 14651 30496 14971 31520
rect 14651 30432 14659 30496
rect 14723 30432 14739 30496
rect 14803 30432 14819 30496
rect 14883 30432 14899 30496
rect 14963 30432 14971 30496
rect 14651 29408 14971 30432
rect 14651 29344 14659 29408
rect 14723 29344 14739 29408
rect 14803 29344 14819 29408
rect 14883 29344 14899 29408
rect 14963 29344 14971 29408
rect 14651 28320 14971 29344
rect 14651 28256 14659 28320
rect 14723 28256 14739 28320
rect 14803 28256 14819 28320
rect 14883 28256 14899 28320
rect 14963 28256 14971 28320
rect 14651 27232 14971 28256
rect 14651 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14971 27232
rect 14651 26144 14971 27168
rect 14651 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14971 26144
rect 14651 25056 14971 26080
rect 14651 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14971 25056
rect 14651 23968 14971 24992
rect 14651 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14971 23968
rect 14651 22880 14971 23904
rect 14651 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14971 22880
rect 14651 21792 14971 22816
rect 14651 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14971 21792
rect 14651 20704 14971 21728
rect 14651 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14971 20704
rect 14651 19616 14971 20640
rect 14651 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14971 19616
rect 14651 18528 14971 19552
rect 14651 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14971 18528
rect 14651 17440 14971 18464
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__conb_1  analog_io_control_1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  analog_io_control_2
timestamp 1688980957
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  analog_io_control_3
timestamp 1688980957
transform -1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  analog_io_control_4
timestamp 1688980957
transform -1 0 14536 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  analog_io_control_5
timestamp 1688980957
transform -1 0 14536 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  analog_io_control_6
timestamp 1688980957
transform -1 0 14536 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_141 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_137 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_145
timestamp 1688980957
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_145
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_145
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_145
timestamp 1688980957
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1688980957
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_145
timestamp 1688980957
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 1688980957
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_145
timestamp 1688980957
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_145
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_145
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_145
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_145
timestamp 1688980957
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1688980957
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_145
timestamp 1688980957
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_145
timestamp 1688980957
transform 1 0 14444 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_145
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_145
timestamp 1688980957
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_145
timestamp 1688980957
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_145
timestamp 1688980957
transform 1 0 14444 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_145
timestamp 1688980957
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_145
timestamp 1688980957
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_145
timestamp 1688980957
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_145
timestamp 1688980957
transform 1 0 14444 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_145
timestamp 1688980957
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_145
timestamp 1688980957
transform 1 0 14444 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_145
timestamp 1688980957
transform 1 0 14444 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_145
timestamp 1688980957
transform 1 0 14444 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_145
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_145
timestamp 1688980957
transform 1 0 14444 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_145
timestamp 1688980957
transform 1 0 14444 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_145
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_145
timestamp 1688980957
transform 1 0 14444 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_145
timestamp 1688980957
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_145
timestamp 1688980957
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_145
timestamp 1688980957
transform 1 0 14444 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_145
timestamp 1688980957
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_145
timestamp 1688980957
transform 1 0 14444 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_145
timestamp 1688980957
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_145
timestamp 1688980957
transform 1 0 14444 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_145
timestamp 1688980957
transform 1 0 14444 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_145
timestamp 1688980957
transform 1 0 14444 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_145
timestamp 1688980957
transform 1 0 14444 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_145
timestamp 1688980957
transform 1 0 14444 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_145
timestamp 1688980957
transform 1 0 14444 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_145
timestamp 1688980957
transform 1 0 14444 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_145
timestamp 1688980957
transform 1 0 14444 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_145
timestamp 1688980957
transform 1 0 14444 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_145
timestamp 1688980957
transform 1 0 14444 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_145
timestamp 1688980957
transform 1 0 14444 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_145
timestamp 1688980957
transform 1 0 14444 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_145
timestamp 1688980957
transform 1 0 14444 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_145
timestamp 1688980957
transform 1 0 14444 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_145
timestamp 1688980957
transform 1 0 14444 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_145
timestamp 1688980957
transform 1 0 14444 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_145
timestamp 1688980957
transform 1 0 14444 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_145
timestamp 1688980957
transform 1 0 14444 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_145
timestamp 1688980957
transform 1 0 14444 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_145
timestamp 1688980957
transform 1 0 14444 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_145
timestamp 1688980957
transform 1 0 14444 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_145
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1688980957
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1688980957
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1688980957
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1688980957
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1688980957
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1688980957
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1688980957
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1688980957
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1688980957
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 1688980957
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1688980957
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_137
timestamp 1688980957
transform 1 0 13708 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_145
timestamp 1688980957
transform 1 0 14444 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1688980957
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1688980957
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1688980957
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1688980957
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1688980957
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1688980957
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1688980957
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_141
timestamp 1688980957
transform 1 0 14076 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_145
timestamp 1688980957
transform 1 0 14444 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_29
timestamp 1688980957
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_41
timestamp 1688980957
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_53
timestamp 1688980957
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1688980957
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_81
timestamp 1688980957
transform 1 0 8556 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_85
timestamp 1688980957
transform 1 0 8924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_97
timestamp 1688980957
transform 1 0 10028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_109
timestamp 1688980957
transform 1 0 11132 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1688980957
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79_137
timestamp 1688980957
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_141
timestamp 1688980957
transform 1 0 14076 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_145
timestamp 1688980957
transform 1 0 14444 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 14812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 14812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 14812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 14812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 14812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 14812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 14812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 14812 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 14812 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 14812 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 14812 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 14812 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 14812 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 14812 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 14812 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 14812 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 14812 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 14812 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 14812 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 14812 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 14812 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 14812 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 14812 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 14812 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 14812 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 14812 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 14812 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 14812 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 3680 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 8832 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 13984 0 -1 45696
box -38 -48 130 592
<< labels >>
flabel metal3 s 15200 4088 16000 4208 0 FreeSans 480 0 0 0 io_oeb[0]
port 0 nsew signal tristate
flabel metal3 s 15200 11976 16000 12096 0 FreeSans 480 0 0 0 io_oeb[1]
port 1 nsew signal tristate
flabel metal3 s 15200 19864 16000 19984 0 FreeSans 480 0 0 0 io_oeb[2]
port 2 nsew signal tristate
flabel metal3 s 15200 27752 16000 27872 0 FreeSans 480 0 0 0 io_oeb[3]
port 3 nsew signal tristate
flabel metal3 s 15200 35640 16000 35760 0 FreeSans 480 0 0 0 io_oeb[4]
port 4 nsew signal tristate
flabel metal3 s 15200 43528 16000 43648 0 FreeSans 480 0 0 0 io_oeb[5]
port 5 nsew signal tristate
flabel metal4 s 2657 2128 2977 45744 0 FreeSans 1920 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 6084 2128 6404 45744 0 FreeSans 1920 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 9511 2128 9831 45744 0 FreeSans 1920 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 12938 2128 13258 45744 0 FreeSans 1920 90 0 0 vccd1
port 6 nsew power bidirectional
flabel metal4 s 4370 2128 4690 45744 0 FreeSans 1920 90 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 45744 0 FreeSans 1920 90 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 45744 0 FreeSans 1920 90 0 0 vssd1
port 7 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 45744 0 FreeSans 1920 90 0 0 vssd1
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 48000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 578.870 BY 589.590 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 10.240 578.870 10.840 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 354.320 578.870 354.920 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 249.600 578.870 250.200 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 70.080 578.870 70.680 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 85.040 578.870 85.640 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 100.000 578.870 100.600 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 114.960 578.870 115.560 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 129.920 578.870 130.520 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 144.880 578.870 145.480 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 159.840 578.870 160.440 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 174.800 578.870 175.400 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 189.760 578.870 190.360 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 204.720 578.870 205.320 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 219.680 578.870 220.280 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 234.640 578.870 235.240 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 264.560 578.870 265.160 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 279.520 578.870 280.120 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 294.480 578.870 295.080 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 309.440 578.870 310.040 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 324.400 578.870 325.000 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 339.360 578.870 339.960 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 369.280 578.870 369.880 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 384.240 578.870 384.840 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 399.200 578.870 399.800 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 414.160 578.870 414.760 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 429.120 578.870 429.720 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 444.080 578.870 444.680 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 459.040 578.870 459.640 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 474.000 578.870 474.600 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 488.960 578.870 489.560 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 503.920 578.870 504.520 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 518.880 578.870 519.480 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 533.840 578.870 534.440 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 548.800 578.870 549.400 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 563.760 578.870 564.360 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 578.720 578.870 579.320 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 25.200 578.870 25.800 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 40.160 578.870 40.760 ;
    END
  END i_reg_mosi
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 574.870 55.120 578.870 55.720 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END i_reset_lock_b
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 585.590 44.070 589.590 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 585.590 32.110 589.590 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 585.590 20.150 589.590 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 585.590 8.190 589.590 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 585.590 115.830 589.590 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 585.590 103.870 589.590 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 585.590 91.910 589.590 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 585.590 79.950 589.590 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 585.590 67.990 589.590 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 585.590 56.030 589.590 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 585.590 187.590 589.590 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 585.590 163.670 589.590 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 585.590 151.710 589.590 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 585.590 139.750 589.590 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 585.590 127.790 589.590 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 585.590 175.630 589.590 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 585.590 570.310 589.590 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 585.590 450.710 589.590 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 585.590 438.750 589.590 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 585.590 426.790 589.590 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 585.590 414.830 589.590 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 585.590 402.870 589.590 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 585.590 390.910 589.590 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 585.590 558.350 589.590 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 585.590 546.390 589.590 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 585.590 534.430 589.590 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 585.590 522.470 589.590 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 585.590 510.510 589.590 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 585.590 498.550 589.590 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 585.590 486.590 589.590 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 585.590 474.630 589.590 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 585.590 462.670 589.590 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 576.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 576.880 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 585.590 378.950 589.590 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 585.590 259.350 589.590 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 585.590 247.390 589.590 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 585.590 235.430 589.590 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 585.590 223.470 589.590 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 585.590 211.510 589.590 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 585.590 199.550 589.590 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 585.590 366.990 589.590 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 585.590 355.030 589.590 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 585.590 343.070 589.590 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 585.590 331.110 589.590 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 585.590 319.150 589.590 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 585.590 307.190 589.590 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 585.590 295.230 589.590 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 585.590 283.270 589.590 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 585.590 271.310 589.590 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 572.505 573.350 575.335 ;
        RECT 5.330 567.065 573.350 569.895 ;
        RECT 5.330 561.625 573.350 564.455 ;
        RECT 5.330 556.185 573.350 559.015 ;
        RECT 5.330 550.745 573.350 553.575 ;
        RECT 5.330 545.305 573.350 548.135 ;
        RECT 5.330 539.865 573.350 542.695 ;
        RECT 5.330 534.425 573.350 537.255 ;
        RECT 5.330 528.985 573.350 531.815 ;
        RECT 5.330 523.545 573.350 526.375 ;
        RECT 5.330 518.105 573.350 520.935 ;
        RECT 5.330 512.665 573.350 515.495 ;
        RECT 5.330 507.225 573.350 510.055 ;
        RECT 5.330 501.785 573.350 504.615 ;
        RECT 5.330 496.345 573.350 499.175 ;
        RECT 5.330 490.905 573.350 493.735 ;
        RECT 5.330 485.465 573.350 488.295 ;
        RECT 5.330 480.025 573.350 482.855 ;
        RECT 5.330 474.585 573.350 477.415 ;
        RECT 5.330 469.145 573.350 471.975 ;
        RECT 5.330 463.705 573.350 466.535 ;
        RECT 5.330 458.265 573.350 461.095 ;
        RECT 5.330 452.825 573.350 455.655 ;
        RECT 5.330 447.385 573.350 450.215 ;
        RECT 5.330 441.945 573.350 444.775 ;
        RECT 5.330 436.505 573.350 439.335 ;
        RECT 5.330 431.065 573.350 433.895 ;
        RECT 5.330 425.625 573.350 428.455 ;
        RECT 5.330 420.185 573.350 423.015 ;
        RECT 5.330 414.745 573.350 417.575 ;
        RECT 5.330 409.305 573.350 412.135 ;
        RECT 5.330 403.865 573.350 406.695 ;
        RECT 5.330 398.425 573.350 401.255 ;
        RECT 5.330 392.985 573.350 395.815 ;
        RECT 5.330 387.545 573.350 390.375 ;
        RECT 5.330 382.105 573.350 384.935 ;
        RECT 5.330 376.665 573.350 379.495 ;
        RECT 5.330 371.225 573.350 374.055 ;
        RECT 5.330 365.785 573.350 368.615 ;
        RECT 5.330 360.345 573.350 363.175 ;
        RECT 5.330 354.905 573.350 357.735 ;
        RECT 5.330 349.465 573.350 352.295 ;
        RECT 5.330 344.025 573.350 346.855 ;
        RECT 5.330 338.585 573.350 341.415 ;
        RECT 5.330 333.145 573.350 335.975 ;
        RECT 5.330 327.705 573.350 330.535 ;
        RECT 5.330 322.265 573.350 325.095 ;
        RECT 5.330 316.825 573.350 319.655 ;
        RECT 5.330 311.385 573.350 314.215 ;
        RECT 5.330 305.945 573.350 308.775 ;
        RECT 5.330 300.505 573.350 303.335 ;
        RECT 5.330 295.065 573.350 297.895 ;
        RECT 5.330 289.625 573.350 292.455 ;
        RECT 5.330 284.185 573.350 287.015 ;
        RECT 5.330 278.745 573.350 281.575 ;
        RECT 5.330 273.305 573.350 276.135 ;
        RECT 5.330 267.865 573.350 270.695 ;
        RECT 5.330 262.425 573.350 265.255 ;
        RECT 5.330 256.985 573.350 259.815 ;
        RECT 5.330 251.545 573.350 254.375 ;
        RECT 5.330 246.105 573.350 248.935 ;
        RECT 5.330 240.665 573.350 243.495 ;
        RECT 5.330 235.225 573.350 238.055 ;
        RECT 5.330 229.785 573.350 232.615 ;
        RECT 5.330 224.345 573.350 227.175 ;
        RECT 5.330 218.905 573.350 221.735 ;
        RECT 5.330 213.465 573.350 216.295 ;
        RECT 5.330 208.025 573.350 210.855 ;
        RECT 5.330 202.585 573.350 205.415 ;
        RECT 5.330 197.145 573.350 199.975 ;
        RECT 5.330 191.705 573.350 194.535 ;
        RECT 5.330 186.265 573.350 189.095 ;
        RECT 5.330 180.825 573.350 183.655 ;
        RECT 5.330 175.385 573.350 178.215 ;
        RECT 5.330 169.945 573.350 172.775 ;
        RECT 5.330 164.505 573.350 167.335 ;
        RECT 5.330 159.065 573.350 161.895 ;
        RECT 5.330 153.625 573.350 156.455 ;
        RECT 5.330 148.185 573.350 151.015 ;
        RECT 5.330 142.745 573.350 145.575 ;
        RECT 5.330 137.305 573.350 140.135 ;
        RECT 5.330 131.865 573.350 134.695 ;
        RECT 5.330 126.425 573.350 129.255 ;
        RECT 5.330 120.985 573.350 123.815 ;
        RECT 5.330 115.545 573.350 118.375 ;
        RECT 5.330 110.105 573.350 112.935 ;
        RECT 5.330 104.665 573.350 107.495 ;
        RECT 5.330 99.225 573.350 102.055 ;
        RECT 5.330 93.785 573.350 96.615 ;
        RECT 5.330 88.345 573.350 91.175 ;
        RECT 5.330 82.905 573.350 85.735 ;
        RECT 5.330 77.465 573.350 80.295 ;
        RECT 5.330 72.025 573.350 74.855 ;
        RECT 5.330 66.585 573.350 69.415 ;
        RECT 5.330 61.145 573.350 63.975 ;
        RECT 5.330 55.705 573.350 58.535 ;
        RECT 5.330 50.265 573.350 53.095 ;
        RECT 5.330 44.825 573.350 47.655 ;
        RECT 5.330 39.385 573.350 42.215 ;
        RECT 5.330 33.945 573.350 36.775 ;
        RECT 5.330 28.505 573.350 31.335 ;
        RECT 5.330 23.065 573.350 25.895 ;
        RECT 5.330 17.625 573.350 20.455 ;
        RECT 5.330 12.185 573.350 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 573.160 576.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 573.460 577.280 ;
      LAYER met2 ;
        RECT 8.470 585.310 19.590 585.590 ;
        RECT 20.430 585.310 31.550 585.590 ;
        RECT 32.390 585.310 43.510 585.590 ;
        RECT 44.350 585.310 55.470 585.590 ;
        RECT 56.310 585.310 67.430 585.590 ;
        RECT 68.270 585.310 79.390 585.590 ;
        RECT 80.230 585.310 91.350 585.590 ;
        RECT 92.190 585.310 103.310 585.590 ;
        RECT 104.150 585.310 115.270 585.590 ;
        RECT 116.110 585.310 127.230 585.590 ;
        RECT 128.070 585.310 139.190 585.590 ;
        RECT 140.030 585.310 151.150 585.590 ;
        RECT 151.990 585.310 163.110 585.590 ;
        RECT 163.950 585.310 175.070 585.590 ;
        RECT 175.910 585.310 187.030 585.590 ;
        RECT 187.870 585.310 198.990 585.590 ;
        RECT 199.830 585.310 210.950 585.590 ;
        RECT 211.790 585.310 222.910 585.590 ;
        RECT 223.750 585.310 234.870 585.590 ;
        RECT 235.710 585.310 246.830 585.590 ;
        RECT 247.670 585.310 258.790 585.590 ;
        RECT 259.630 585.310 270.750 585.590 ;
        RECT 271.590 585.310 282.710 585.590 ;
        RECT 283.550 585.310 294.670 585.590 ;
        RECT 295.510 585.310 306.630 585.590 ;
        RECT 307.470 585.310 318.590 585.590 ;
        RECT 319.430 585.310 330.550 585.590 ;
        RECT 331.390 585.310 342.510 585.590 ;
        RECT 343.350 585.310 354.470 585.590 ;
        RECT 355.310 585.310 366.430 585.590 ;
        RECT 367.270 585.310 378.390 585.590 ;
        RECT 379.230 585.310 390.350 585.590 ;
        RECT 391.190 585.310 402.310 585.590 ;
        RECT 403.150 585.310 414.270 585.590 ;
        RECT 415.110 585.310 426.230 585.590 ;
        RECT 427.070 585.310 438.190 585.590 ;
        RECT 439.030 585.310 450.150 585.590 ;
        RECT 450.990 585.310 462.110 585.590 ;
        RECT 462.950 585.310 474.070 585.590 ;
        RECT 474.910 585.310 486.030 585.590 ;
        RECT 486.870 585.310 497.990 585.590 ;
        RECT 498.830 585.310 509.950 585.590 ;
        RECT 510.790 585.310 521.910 585.590 ;
        RECT 522.750 585.310 533.870 585.590 ;
        RECT 534.710 585.310 545.830 585.590 ;
        RECT 546.670 585.310 557.790 585.590 ;
        RECT 558.630 585.310 569.750 585.590 ;
        RECT 570.590 585.310 571.680 585.590 ;
        RECT 7.920 4.280 571.680 585.310 ;
        RECT 7.920 4.000 8.090 4.280 ;
        RECT 8.930 4.000 23.270 4.280 ;
        RECT 24.110 4.000 38.450 4.280 ;
        RECT 39.290 4.000 53.630 4.280 ;
        RECT 54.470 4.000 68.810 4.280 ;
        RECT 69.650 4.000 83.990 4.280 ;
        RECT 84.830 4.000 99.170 4.280 ;
        RECT 100.010 4.000 114.350 4.280 ;
        RECT 115.190 4.000 129.530 4.280 ;
        RECT 130.370 4.000 144.710 4.280 ;
        RECT 145.550 4.000 159.890 4.280 ;
        RECT 160.730 4.000 175.070 4.280 ;
        RECT 175.910 4.000 190.250 4.280 ;
        RECT 191.090 4.000 205.430 4.280 ;
        RECT 206.270 4.000 220.610 4.280 ;
        RECT 221.450 4.000 235.790 4.280 ;
        RECT 236.630 4.000 250.970 4.280 ;
        RECT 251.810 4.000 266.150 4.280 ;
        RECT 266.990 4.000 281.330 4.280 ;
        RECT 282.170 4.000 296.510 4.280 ;
        RECT 297.350 4.000 311.690 4.280 ;
        RECT 312.530 4.000 326.870 4.280 ;
        RECT 327.710 4.000 342.050 4.280 ;
        RECT 342.890 4.000 357.230 4.280 ;
        RECT 358.070 4.000 372.410 4.280 ;
        RECT 373.250 4.000 387.590 4.280 ;
        RECT 388.430 4.000 402.770 4.280 ;
        RECT 403.610 4.000 417.950 4.280 ;
        RECT 418.790 4.000 433.130 4.280 ;
        RECT 433.970 4.000 448.310 4.280 ;
        RECT 449.150 4.000 463.490 4.280 ;
        RECT 464.330 4.000 478.670 4.280 ;
        RECT 479.510 4.000 493.850 4.280 ;
        RECT 494.690 4.000 509.030 4.280 ;
        RECT 509.870 4.000 524.210 4.280 ;
        RECT 525.050 4.000 539.390 4.280 ;
        RECT 540.230 4.000 554.570 4.280 ;
        RECT 555.410 4.000 569.750 4.280 ;
        RECT 570.590 4.000 571.680 4.280 ;
      LAYER met3 ;
        RECT 21.050 578.320 574.470 579.185 ;
        RECT 21.050 564.760 574.870 578.320 ;
        RECT 21.050 563.360 574.470 564.760 ;
        RECT 21.050 549.800 574.870 563.360 ;
        RECT 21.050 548.400 574.470 549.800 ;
        RECT 21.050 534.840 574.870 548.400 ;
        RECT 21.050 533.440 574.470 534.840 ;
        RECT 21.050 519.880 574.870 533.440 ;
        RECT 21.050 518.480 574.470 519.880 ;
        RECT 21.050 504.920 574.870 518.480 ;
        RECT 21.050 503.520 574.470 504.920 ;
        RECT 21.050 489.960 574.870 503.520 ;
        RECT 21.050 488.560 574.470 489.960 ;
        RECT 21.050 475.000 574.870 488.560 ;
        RECT 21.050 473.600 574.470 475.000 ;
        RECT 21.050 460.040 574.870 473.600 ;
        RECT 21.050 458.640 574.470 460.040 ;
        RECT 21.050 445.080 574.870 458.640 ;
        RECT 21.050 443.680 574.470 445.080 ;
        RECT 21.050 430.120 574.870 443.680 ;
        RECT 21.050 428.720 574.470 430.120 ;
        RECT 21.050 415.160 574.870 428.720 ;
        RECT 21.050 413.760 574.470 415.160 ;
        RECT 21.050 400.200 574.870 413.760 ;
        RECT 21.050 398.800 574.470 400.200 ;
        RECT 21.050 385.240 574.870 398.800 ;
        RECT 21.050 383.840 574.470 385.240 ;
        RECT 21.050 370.280 574.870 383.840 ;
        RECT 21.050 368.880 574.470 370.280 ;
        RECT 21.050 355.320 574.870 368.880 ;
        RECT 21.050 353.920 574.470 355.320 ;
        RECT 21.050 340.360 574.870 353.920 ;
        RECT 21.050 338.960 574.470 340.360 ;
        RECT 21.050 325.400 574.870 338.960 ;
        RECT 21.050 324.000 574.470 325.400 ;
        RECT 21.050 310.440 574.870 324.000 ;
        RECT 21.050 309.040 574.470 310.440 ;
        RECT 21.050 295.480 574.870 309.040 ;
        RECT 21.050 294.080 574.470 295.480 ;
        RECT 21.050 280.520 574.870 294.080 ;
        RECT 21.050 279.120 574.470 280.520 ;
        RECT 21.050 265.560 574.870 279.120 ;
        RECT 21.050 264.160 574.470 265.560 ;
        RECT 21.050 250.600 574.870 264.160 ;
        RECT 21.050 249.200 574.470 250.600 ;
        RECT 21.050 235.640 574.870 249.200 ;
        RECT 21.050 234.240 574.470 235.640 ;
        RECT 21.050 220.680 574.870 234.240 ;
        RECT 21.050 219.280 574.470 220.680 ;
        RECT 21.050 205.720 574.870 219.280 ;
        RECT 21.050 204.320 574.470 205.720 ;
        RECT 21.050 190.760 574.870 204.320 ;
        RECT 21.050 189.360 574.470 190.760 ;
        RECT 21.050 175.800 574.870 189.360 ;
        RECT 21.050 174.400 574.470 175.800 ;
        RECT 21.050 160.840 574.870 174.400 ;
        RECT 21.050 159.440 574.470 160.840 ;
        RECT 21.050 145.880 574.870 159.440 ;
        RECT 21.050 144.480 574.470 145.880 ;
        RECT 21.050 130.920 574.870 144.480 ;
        RECT 21.050 129.520 574.470 130.920 ;
        RECT 21.050 115.960 574.870 129.520 ;
        RECT 21.050 114.560 574.470 115.960 ;
        RECT 21.050 101.000 574.870 114.560 ;
        RECT 21.050 99.600 574.470 101.000 ;
        RECT 21.050 86.040 574.870 99.600 ;
        RECT 21.050 84.640 574.470 86.040 ;
        RECT 21.050 71.080 574.870 84.640 ;
        RECT 21.050 69.680 574.470 71.080 ;
        RECT 21.050 56.120 574.870 69.680 ;
        RECT 21.050 54.720 574.470 56.120 ;
        RECT 21.050 41.160 574.870 54.720 ;
        RECT 21.050 39.760 574.470 41.160 ;
        RECT 21.050 26.200 574.870 39.760 ;
        RECT 21.050 24.800 574.470 26.200 ;
        RECT 21.050 11.240 574.870 24.800 ;
        RECT 21.050 9.840 574.470 11.240 ;
        RECT 21.050 9.695 574.870 9.840 ;
      LAYER met4 ;
        RECT 78.495 10.240 97.440 566.945 ;
        RECT 99.840 10.240 174.240 566.945 ;
        RECT 176.640 10.240 251.040 566.945 ;
        RECT 253.440 10.240 327.840 566.945 ;
        RECT 330.240 10.240 404.640 566.945 ;
        RECT 407.040 10.240 481.440 566.945 ;
        RECT 483.840 10.240 492.825 566.945 ;
        RECT 78.495 9.695 492.825 10.240 ;
  END
END top_ew_algofoogle
END LIBRARY

